* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : nand2                                        *
* Netlisted  : Wed Dec  3 20:57:04 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764817018881                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764817018881 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764817018881

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764817018883                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764817018883 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764817018883

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764817018880                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764817018880 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764817018880

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764817018881                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764817018881 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_764817018881

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand2                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand2 3 4 2 6 5
** N=6 EP=5 FDC=8
X0 1 M2_M1_CDNS_764817018881 $T=230 -2010 0 0 $X=150 $Y=-2260
X1 2 M2_M1_CDNS_764817018881 $T=640 860 0 0 $X=560 $Y=610
X2 1 M2_M1_CDNS_764817018881 $T=1050 -2010 0 0 $X=970 $Y=-2260
X3 1 M2_M1_CDNS_764817018881 $T=1530 -2010 0 0 $X=1450 $Y=-2260
X4 2 M2_M1_CDNS_764817018881 $T=1940 860 0 0 $X=1860 $Y=610
X5 1 M2_M1_CDNS_764817018881 $T=2350 -2010 0 0 $X=2270 $Y=-2260
X6 3 M1_PO_CDNS_764817018883 $T=290 -430 0 0 $X=190 $Y=-790
X7 4 M1_PO_CDNS_764817018883 $T=1590 -730 0 0 $X=1490 $Y=-1090
X8 1 1 2 3 5 nmos1v_CDNS_764817018880 $T=390 -2730 0 0 $X=-30 $Y=-2930
X9 1 1 5 4 5 nmos1v_CDNS_764817018880 $T=1690 -2730 0 0 $X=1270 $Y=-2930
X10 2 6 6 3 5 6 pmos1v_CDNS_764817018881 $T=390 140 0 0 $X=-30 $Y=-60
X11 2 6 6 4 5 6 pmos1v_CDNS_764817018881 $T=1690 140 0 0 $X=1270 $Y=-60
M0 2 3 6 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=390 $Y=140 $dt=1
M1 6 3 2 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.4011 scb=0.0195321 scc=0.00239618 $X=800 $Y=140 $dt=1
M2 2 4 6 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.4011 scb=0.0195321 scc=0.00239618 $X=1690 $Y=140 $dt=1
M3 6 4 2 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2100 $Y=140 $dt=1
.ends nand2
