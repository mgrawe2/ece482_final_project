* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : full_adder                                   *
* Netlisted  : Sun Nov 30 12:11:44 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764526298900                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764526298900 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764526298900

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764526298901                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764526298901 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764526298901

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764526298902                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764526298902 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764526298902

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764526298905                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764526298905 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764526298905

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764526298907                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764526298907 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764526298907

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764526298908                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764526298908 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764526298908

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764526298909                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764526298909 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764526298909

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7645262989010                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7645262989010 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7645262989010

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7645262989011                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7645262989011 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7645262989011

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7645262989012                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7645262989012 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7645262989012

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7645262989013                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7645262989013 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7645262989013

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7645262989014                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7645262989014 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7645262989014

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_7645262989015                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_7645262989015 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_7645262989015

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_7645262989016                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_7645262989016 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_7645262989016

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_7645262989017                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_7645262989017 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_7645262989017

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_7645262989018                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_7645262989018 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_7645262989018

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764526298900                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764526298900 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 3 1 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=7.55e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=0 $Y=0 $dt=1
M1 4 6 2 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=5.5e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=410 $Y=0 $dt=1
M2 5 7 4 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=3.45e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=820 $Y=0 $dt=1
M3 8 9 5 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=7.55e-07 sb=1.4e-07 sca=30.82 scb=0.02528 scc=0.00362484 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_764526298900

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764526298901                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764526298901 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_764526298901

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764526298902                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764526298902 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_764526298902

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764526298903                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764526298903 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764526298903

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
X0 4 3 1 nmos1v_CDNS_764526298902 $T=-50 -540 0 0 $X=-470 $Y=-740
X1 2 3 1 4 2 pmos1v_CDNS_764526298903 $T=-50 460 0 0 $X=-470 $Y=260
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764526298904                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764526298904 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=0 $Y=0 $dt=1
M1 3 1 2 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=410 $Y=0 $dt=1
.ends pmos1v_CDNS_764526298904

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764526298905                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764526298905 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=0 $Y=0 $dt=0
M1 3 1 2 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764526298905

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=5
X0 5 M1_PO_CDNS_764526298900 $T=850 -1090 0 0 $X=750 $Y=-1450
X1 1 M1_PO_CDNS_764526298900 $T=850 2390 0 0 $X=750 $Y=2030
X2 4 M1_PO_CDNS_764526298900 $T=1260 650 0 0 $X=1160 $Y=290
X3 4 M2_M1_CDNS_764526298908 $T=360 650 0 0 $X=280 $Y=240
X4 4 M2_M1_CDNS_764526298908 $T=1260 650 0 0 $X=1180 $Y=240
X5 1 2 5 3 inv $T=-790 -50 0 0 $X=-1590 $Y=-1230
X6 4 6 1 3 2 pmos1v_CDNS_764526298904 $T=660 1350 0 0 $X=240 $Y=1150
X7 4 6 5 3 nmos1v_CDNS_764526298905 $T=660 -340 0 0 $X=240 $Y=-540
M0 5 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.6083 scb=0.0129915 scc=0.000573075 $X=-840 $Y=-590 $dt=0
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 4 8 1 10 5 7 9
** N=15 EP=7 FDC=22
X0 1 M1_PO_CDNS_764526298900 $T=790 -2720 0 0 $X=690 $Y=-3080
X1 2 M1_PO_CDNS_764526298900 $T=1490 -1360 0 0 $X=1390 $Y=-1720
X2 3 M1_PO_CDNS_764526298900 $T=1490 -160 0 0 $X=1390 $Y=-520
X3 3 M1_PO_CDNS_764526298900 $T=1900 -1360 0 0 $X=1800 $Y=-1720
X4 2 M1_PO_CDNS_764526298900 $T=1900 -160 0 0 $X=1800 $Y=-520
X5 4 M1_PO_CDNS_764526298900 $T=2310 -2720 0 0 $X=2210 $Y=-3080
X6 2 M2_M1_CDNS_764526298901 $T=-4410 -500 0 0 $X=-4490 $Y=-770
X7 5 M2_M1_CDNS_764526298901 $T=-610 -540 0 0 $X=-690 $Y=-810
X8 3 M2_M1_CDNS_764526298901 $T=-540 -2000 0 0 $X=-620 $Y=-2270
X9 6 M2_M1_CDNS_764526298901 $T=590 -90 0 0 $X=510 $Y=-360
X10 1 M2_M1_CDNS_764526298901 $T=790 -2710 0 0 $X=710 $Y=-2980
X11 2 M2_M1_CDNS_764526298901 $T=1490 -1390 0 0 $X=1410 $Y=-1660
X12 3 M2_M1_CDNS_764526298901 $T=1900 -1360 0 0 $X=1820 $Y=-1630
X13 2 M2_M1_CDNS_764526298901 $T=1900 -160 0 0 $X=1820 $Y=-430
X14 4 M2_M1_CDNS_764526298901 $T=2320 -2720 0 0 $X=2240 $Y=-2990
X15 6 M2_M1_CDNS_764526298901 $T=2510 -70 0 0 $X=2430 $Y=-340
X16 2 M3_M2_CDNS_764526298902 $T=-4410 -500 0 0 $X=-4490 $Y=-770
X17 5 M3_M2_CDNS_764526298902 $T=-610 -540 0 0 $X=-690 $Y=-810
X18 3 M3_M2_CDNS_764526298902 $T=-540 -2000 0 0 $X=-620 $Y=-2270
X19 6 M3_M2_CDNS_764526298902 $T=590 -90 0 0 $X=510 $Y=-360
X20 1 M3_M2_CDNS_764526298902 $T=790 -2710 0 0 $X=710 $Y=-2980
X21 3 M3_M2_CDNS_764526298902 $T=1900 -1360 0 0 $X=1820 $Y=-1630
X22 6 M3_M2_CDNS_764526298902 $T=2510 -70 0 0 $X=2430 $Y=-340
X23 7 M2_M1_CDNS_764526298905 $T=-6190 480 0 0 $X=-6410 $Y=350
X24 2 M2_M1_CDNS_764526298905 $T=-2450 -890 0 0 $X=-2670 $Y=-1020
X25 7 M2_M1_CDNS_764526298905 $T=-2390 480 0 0 $X=-2610 $Y=350
X26 7 M2_M1_CDNS_764526298905 $T=1530 1390 0 0 $X=1310 $Y=1260
X27 8 M3_M2_CDNS_764526298907 $T=-6990 -3990 0 0 $X=-7070 $Y=-4400
X28 4 M3_M2_CDNS_764526298907 $T=-4300 -3990 0 0 $X=-4380 $Y=-4400
X29 1 M3_M2_CDNS_764526298907 $T=-1030 -260 0 0 $X=-1110 $Y=-670
X30 5 M3_M2_CDNS_764526298907 $T=-600 2400 0 0 $X=-680 $Y=1990
X31 8 M2_M1_CDNS_764526298908 $T=-6990 -3990 0 0 $X=-7070 $Y=-4400
X32 4 M2_M1_CDNS_764526298908 $T=-4300 -3990 0 0 $X=-4380 $Y=-4400
X33 5 M2_M1_CDNS_764526298908 $T=-600 2400 0 0 $X=-680 $Y=1990
X34 1 M3_M2_CDNS_764526298909 $T=-7660 -2700 0 0 $X=-8020 $Y=-2830
X35 9 M3_M2_CDNS_764526298909 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X36 7 M3_M2_CDNS_764526298909 $T=3220 2330 0 0 $X=2860 $Y=2200
X37 10 M3_M2_CDNS_764526298909 $T=4650 0 0 0 $X=4290 $Y=-130
X38 1 M2_M1_CDNS_7645262989010 $T=-7660 -2700 0 0 $X=-8020 $Y=-2830
X39 9 M2_M1_CDNS_7645262989010 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X40 7 M2_M1_CDNS_7645262989010 $T=3220 2330 0 0 $X=2860 $Y=2200
X41 10 M2_M1_CDNS_7645262989010 $T=4650 0 0 0 $X=4290 $Y=-130
X42 9 M4_M3_CDNS_7645262989011 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X43 7 M4_M3_CDNS_7645262989011 $T=3220 2330 0 0 $X=2860 $Y=2200
X44 9 M5_M4_CDNS_7645262989012 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X45 7 M5_M4_CDNS_7645262989012 $T=3220 2330 0 0 $X=2860 $Y=2200
X46 9 M6_M5_CDNS_7645262989013 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X47 7 M6_M5_CDNS_7645262989013 $T=3220 2330 0 0 $X=2860 $Y=2200
X48 9 M7_M6_CDNS_7645262989014 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X49 7 M7_M6_CDNS_7645262989014 $T=3220 2330 0 0 $X=2860 $Y=2200
X50 9 M8_M7_CDNS_7645262989015 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X51 7 M8_M7_CDNS_7645262989015 $T=3220 2330 0 0 $X=2860 $Y=2200
X52 9 M9_M8_CDNS_7645262989016 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X53 7 M9_M8_CDNS_7645262989016 $T=3220 2330 0 0 $X=2860 $Y=2200
X54 9 M10_M9_CDNS_7645262989017 $T=1590 -4010 0 0 $X=630 $Y=-4290
X55 7 M10_M9_CDNS_7645262989017 $T=3240 2340 0 0 $X=2280 $Y=2060
X56 9 M11_M10_CDNS_7645262989018 $T=1590 -4010 0 0 $X=630 $Y=-4290
X57 7 M11_M10_CDNS_7645262989018 $T=3240 2340 0 0 $X=2280 $Y=2060
X58 6 11 1 7 12 3 2 6 4 9
+ 7 pmos1v_CDNS_764526298900 $T=890 400 0 0 $X=470 $Y=200
X59 6 13 1 9 14 2 3 6 4 nmos1v_CDNS_764526298901 $T=890 -2160 0 0 $X=470 $Y=-2360
X60 6 7 10 9 inv $T=3440 20 0 0 $X=2640 $Y=-1160
X61 8 7 9 4 15 2 xor $T=-5190 -910 0 0 $X=-7060 $Y=-2360
X62 2 7 9 1 3 5 xor $T=-1390 -910 0 0 $X=-3260 $Y=-2360
M0 10 6 9 9 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=15.2291 scb=0.0163495 scc=0.00102074 $X=3390 $Y=-520 $dt=0
M1 15 8 7 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=38.1374 scb=0.0367153 scc=0.003591 $X=-6030 $Y=-500 $dt=1
M2 3 2 7 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=37.8604 scb=0.0362251 scc=0.00357304 $X=-2230 $Y=-500 $dt=1
M3 10 6 7 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=28.8254 scb=0.0308995 scc=0.00229409 $X=3390 $Y=480 $dt=1
.ends full_adder
