* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : c2mos                                        *
* Netlisted  : Sun Dec  7 19:23:32 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765157006930                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765157006930 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765157006930

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765157006931                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765157006931 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765157006931

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765157006932                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765157006932 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765157006932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765157006930                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765157006930 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765157006930

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765157006931                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765157006931 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765157006931

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765157006932                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765157006932 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765157006932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: c2mos                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt c2mos 1 4 10 5 6 7
** N=12 EP=6 FDC=11
X0 1 M2_M1_CDNS_765157006930 $T=480 1970 0 90 $X=350 $Y=1890
X1 2 M2_M1_CDNS_765157006930 $T=1070 1420 0 90 $X=940 $Y=1340
X2 1 M2_M1_CDNS_765157006930 $T=3650 1970 0 90 $X=3520 $Y=1890
X3 2 M2_M1_CDNS_765157006930 $T=3660 1420 0 90 $X=3530 $Y=1340
X4 3 M2_M1_CDNS_765157006930 $T=4060 1720 0 90 $X=3930 $Y=1640
X5 3 M2_M1_CDNS_765157006930 $T=5220 1720 0 90 $X=5090 $Y=1640
X6 1 M2_M1_CDNS_765157006930 $T=5960 2040 0 90 $X=5830 $Y=1960
X7 2 M2_M1_CDNS_765157006930 $T=6620 1970 0 90 $X=6490 $Y=1890
X8 1 M1_PO_CDNS_765157006931 $T=3660 1980 0 90 $X=3540 $Y=1880
X9 2 M1_PO_CDNS_765157006931 $T=3670 1420 0 90 $X=3550 $Y=1320
X10 3 M1_PO_CDNS_765157006931 $T=5210 1720 0 90 $X=5090 $Y=1620
X11 2 M1_PO_CDNS_765157006931 $T=6630 1980 0 90 $X=6510 $Y=1880
X12 1 M1_PO_CDNS_765157006931 $T=6660 1400 0 90 $X=6540 $Y=1300
X13 1 M1_PO_CDNS_765157006932 $T=530 1970 0 0 $X=310 $Y=1850
X14 4 M1_PO_CDNS_765157006932 $T=2110 1720 0 0 $X=1890 $Y=1600
X15 5 M1_PO_CDNS_765157006932 $T=8090 1590 0 0 $X=7870 $Y=1470
X16 6 2 1 7 6 pmos1v_CDNS_765157006930 $T=750 2360 0 0 $X=330 $Y=2160
X17 6 8 4 7 6 pmos1v_CDNS_765157006930 $T=2240 2360 0 0 $X=1820 $Y=2160
X18 8 3 1 7 6 pmos1v_CDNS_765157006930 $T=3740 2350 0 0 $X=3320 $Y=2150
X19 6 9 3 7 6 pmos1v_CDNS_765157006930 $T=5230 2360 0 0 $X=4810 $Y=2160
X20 9 10 2 7 6 pmos1v_CDNS_765157006930 $T=6720 2340 0 0 $X=6300 $Y=2140
X21 7 1 2 7 nmos1v_CDNS_765157006931 $T=750 650 0 0 $X=330 $Y=450
X22 7 4 11 7 nmos1v_CDNS_765157006931 $T=2240 650 0 0 $X=1820 $Y=450
X23 11 2 3 7 nmos1v_CDNS_765157006931 $T=3750 650 0 0 $X=3330 $Y=450
X24 7 3 12 7 nmos1v_CDNS_765157006931 $T=5230 650 0 0 $X=4810 $Y=450
X25 12 1 10 7 nmos1v_CDNS_765157006931 $T=6720 650 0 0 $X=6300 $Y=450
X26 10 7 5 nmos1v_CDNS_765157006932 $T=8210 170 0 0 $X=7790 $Y=-30
M0 2 1 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.27 scb=0.0231774 scc=0.00199917 $X=750 $Y=2360 $dt=1
M1 8 4 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=2240 $Y=2360 $dt=1
M2 3 1 8 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.7063 scb=0.016025 scc=0.00198503 $X=3740 $Y=2350 $dt=1
M3 9 3 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=5230 $Y=2360 $dt=1
M4 10 2 9 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.6749 scb=0.0214174 scc=0.0021813 $X=6720 $Y=2340 $dt=1
.ends c2mos
