* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mult                                         *
* Netlisted  : Sun Nov 30 19:17:02 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764551816960                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764551816960 S_source_0 D_drain_1 3 S_source_2 D_drain_3 6 7 S_source_4 9 B
** N=11 EP=10 FDC=4
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=7.55e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=0 $Y=0 $dt=1
M1 S_source_2 6 D_drain_1 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=5.5e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=410 $Y=0 $dt=1
M2 D_drain_3 7 S_source_2 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=3.45e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=820 $Y=0 $dt=1
M3 S_source_4 9 D_drain_3 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=7.55e-07 sb=1.4e-07 sca=30.82 scb=0.02528 scc=0.00362484 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_764551816960

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764551816961                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764551816961 S_source_0 D_drain_1 3 S_source_2 D_drain_3 6 7 S_source_4 9
** N=9 EP=9 FDC=4
M0 D_drain_1 3 S_source_0 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 S_source_2 6 D_drain_1 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 D_drain_3 7 S_source_2 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
M3 S_source_4 9 D_drain_3 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_764551816961

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764551816965                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764551816965 S_source_0 D_drain_1 S_source_2 4
** N=4 EP=4 FDC=2
M0 D_drain_1 S_source_2 S_source_0 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=0 $Y=0 $dt=0
M1 S_source_2 S_source_0 D_drain_1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764551816965

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor B VDD VSS 4 B_Bar OUT
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X7 4 OUT B_Bar VSS nmos1v_CDNS_764551816965 $T=660 -340 0 0 $X=240 $Y=-540
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder B Ci VDD VSS A S Co
** N=15 EP=7 FDC=22
X60 10 11 Ci VDD 12 9 8 10 A VDD pmos1v_CDNS_764551816960 $T=890 400 0 0 $X=470 $Y=200
X61 10 13 Ci VSS 14 8 9 10 A nmos1v_CDNS_764551816961 $T=890 -2160 0 0 $X=470 $Y=-2360
X63 B VDD VSS A 15 8 xor $T=-5190 -910 0 0 $X=-7060 $Y=-2360
X64 8 VDD VSS Ci 9 S xor $T=-1390 -910 0 0 $X=-3260 $Y=-2360
M0 15 B VSS VSS g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.6083 scb=0.0129915 scc=0.000573075 $X=-6030 $Y=-1500 $dt=0
M1 9 8 VSS VSS g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.6083 scb=0.0129915 scc=0.000573075 $X=-2230 $Y=-1500 $dt=0
M2 Co 10 VSS VSS g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=15.2291 scb=0.0163495 scc=0.00102074 $X=3390 $Y=-520 $dt=0
M3 15 B VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=38.1374 scb=0.0367153 scc=0.003591 $X=-6030 $Y=-500 $dt=1
M4 8 B A VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-4530 $Y=440 $dt=1
M5 B A 8 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-4120 $Y=440 $dt=1
M6 9 8 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=37.8604 scb=0.0362251 scc=0.00357304 $X=-2230 $Y=-500 $dt=1
M7 S 8 Ci VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-730 $Y=440 $dt=1
M8 8 Ci S VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-320 $Y=440 $dt=1
M9 Co 10 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=28.8254 scb=0.0308995 scc=0.00229409 $X=3390 $Y=480 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764551816967                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764551816967 S_source_0 D_drain_1 3 4 S_source_2 D_drain_3
** N=6 EP=6 FDC=3
M0 D_drain_1 3 S_source_0 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 S_source_2 4 D_drain_1 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 D_drain_3 S_source_0 S_source_2 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
.ends nmos1v_CDNS_764551816967

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 VDD VSS B A OUT 6
*.DEVICECLIMB
** N=7 EP=6 FDC=3
X36 6 7 A B VSS OUT nmos1v_CDNS_764551816967 $T=-460 -1890 0 0 $X=-880 $Y=-2090
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder B VDD VSS A S Co
** N=9 EP=6 FDC=12
X12 B VDD VSS A 7 S xor $T=-2220 70 0 0 $X=-4090 $Y=-1380
X13 VDD VSS B A Co 8 and2 $T=630 630 0 0 $X=-960 $Y=-4060
M0 7 B VSS VSS g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.9282 scb=0.0134361 scc=0.000622896 $X=-3060 $Y=-520 $dt=0
M1 7 B VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=36.6317 scb=0.035909 scc=0.00335548 $X=-3060 $Y=480 $dt=1
M2 S B A VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=-1560 $Y=1420 $dt=1
M3 B A S VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=-1150 $Y=1420 $dt=1
M4 8 A VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=26.2992 scb=0.0240146 scc=0.00255754 $X=170 $Y=1450 $dt=1
M5 VDD B 8 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=28.7383 scb=0.0277231 scc=0.00260208 $X=580 $Y=1450 $dt=1
M6 Co 8 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=39.2498 scb=0.0428135 scc=0.00408073 $X=990 $Y=1450 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mult                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mult A0 A1 A2 A3 B0 B1 B2 B3 P0 P1
+ P2 P3 P4 P5 P6 P7 VDD VSS
** N=142 EP=18 FDC=320
X0 1 2 VDD VSS 5 6 7 full_adder $T=-5100 -5060 0 0 $X=-13120 $Y=-9460
X1 8 9 VDD VSS 10 11 12 full_adder $T=7620 11130 0 0 $X=-400 $Y=6730
X2 13 7 VDD VSS 14 10 15 full_adder $T=8320 -5030 0 0 $X=300 $Y=-9430
X3 16 17 VDD VSS 18 P4 20 full_adder $T=20720 27820 0 0 $X=12700 $Y=23420
X4 21 12 VDD VSS 22 18 23 full_adder $T=21270 11120 0 0 $X=13250 $Y=6720
X5 24 20 VDD VSS 25 P5 27 full_adder $T=34370 27810 0 0 $X=26350 $Y=23410
X6 28 23 VDD VSS 29 25 30 full_adder $T=35050 11120 0 0 $X=27030 $Y=6720
X7 31 27 VDD VSS 30 P6 P7 full_adder $T=48150 27810 0 0 $X=40130 $Y=23410
X8 VDD VSS B0 A0 P0 83 and2 $T=-26670 -21260 0 0 $X=-28260 $Y=-25950
X9 VDD VSS B0 A1 38 84 and2 $T=-22280 -21130 0 0 $X=-23870 $Y=-25820
X10 VDD VSS B1 A0 40 85 and2 $T=-18840 -12210 0 0 $X=-20430 $Y=-16900
X11 VDD VSS B0 A2 5 86 and2 $T=-13020 -21220 0 0 $X=-14610 $Y=-25910
X12 VDD VSS B2 A0 43 87 and2 $T=-12210 3290 0 0 $X=-13800 $Y=-1400
X13 VDD VSS B1 A1 1 88 and2 $T=-10040 -12640 0 0 $X=-11630 $Y=-17330
X14 VDD VSS B2 A1 8 89 and2 $T=400 3630 0 0 $X=-1190 $Y=-1060
X15 VDD VSS B0 A3 14 90 and2 $T=540 -21460 0 0 $X=-1050 $Y=-26150
X16 VDD VSS B3 A0 46 91 and2 $T=890 19980 0 0 $X=-700 $Y=15290
X17 VDD VSS B1 A2 13 92 and2 $T=3520 -12410 0 0 $X=1930 $Y=-17100
X18 VDD VSS B3 A1 16 93 and2 $T=13500 20320 0 0 $X=11910 $Y=15630
X19 VDD VSS B2 A2 21 94 and2 $T=14000 3190 0 0 $X=12410 $Y=-1500
X20 VDD VSS B1 A3 47 95 and2 $T=15640 -12550 0 0 $X=14050 $Y=-17240
X21 VDD VSS B3 A2 24 96 and2 $T=27100 19880 0 0 $X=25510 $Y=15190
X22 VDD VSS B2 A3 28 97 and2 $T=27120 3240 0 0 $X=25530 $Y=-1450
X23 VDD VSS B3 A3 31 98 and2 $T=40220 19930 0 0 $X=38630 $Y=15240
X24 40 VDD VSS 38 P1 2 half_adder $T=-15990 -5900 0 0 $X=-20240 $Y=-9960
X25 43 VDD VSS 6 P2 9 half_adder $T=-7050 9650 0 0 $X=-11300 $Y=5590
X26 46 VDD VSS 11 P3 17 half_adder $T=6050 26340 0 0 $X=1800 $Y=22280
X27 15 VDD VSS 47 22 29 half_adder $T=18470 -5780 0 0 $X=14220 $Y=-9840
M0 83 A0 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-27130 $Y=-20440 $dt=1
M1 VDD B0 83 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-26720 $Y=-20440 $dt=1
M2 P0 83 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-26310 $Y=-20440 $dt=1
M3 84 A1 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-22740 $Y=-20310 $dt=1
M4 VDD B0 84 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-22330 $Y=-20310 $dt=1
M5 38 84 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-21920 $Y=-20310 $dt=1
M6 85 A0 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-19300 $Y=-11390 $dt=1
M7 VDD B1 85 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-18890 $Y=-11390 $dt=1
M8 40 85 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-18480 $Y=-11390 $dt=1
M9 86 A2 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-13480 $Y=-20400 $dt=1
M10 VDD B0 86 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-13070 $Y=-20400 $dt=1
M11 87 A0 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-12670 $Y=4110 $dt=1
M12 5 86 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-12660 $Y=-20400 $dt=1
M13 VDD B2 87 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-12260 $Y=4110 $dt=1
M14 43 87 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-11850 $Y=4110 $dt=1
M15 88 A1 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-10500 $Y=-11820 $dt=1
M16 VDD B1 88 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-10090 $Y=-11820 $dt=1
M17 1 88 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-9680 $Y=-11820 $dt=1
M18 89 A1 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-60 $Y=4450 $dt=1
M19 90 A3 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=80 $Y=-20640 $dt=1
M20 VDD B2 89 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=350 $Y=4450 $dt=1
M21 91 A0 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=430 $Y=20800 $dt=1
M22 VDD B0 90 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=490 $Y=-20640 $dt=1
M23 8 89 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=760 $Y=4450 $dt=1
M24 VDD B3 91 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=840 $Y=20800 $dt=1
M25 14 90 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=900 $Y=-20640 $dt=1
M26 46 91 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=1250 $Y=20800 $dt=1
M27 92 A2 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=3060 $Y=-11590 $dt=1
M28 VDD B1 92 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=3470 $Y=-11590 $dt=1
M29 13 92 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=3880 $Y=-11590 $dt=1
M30 93 A1 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=13040 $Y=21140 $dt=1
M31 VDD B3 93 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=13450 $Y=21140 $dt=1
M32 94 A2 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=13540 $Y=4010 $dt=1
M33 16 93 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=13860 $Y=21140 $dt=1
M34 VDD B2 94 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=13950 $Y=4010 $dt=1
M35 21 94 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=14360 $Y=4010 $dt=1
M36 95 A3 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=15180 $Y=-11730 $dt=1
M37 VDD B1 95 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=15590 $Y=-11730 $dt=1
M38 47 95 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=16000 $Y=-11730 $dt=1
M39 96 A2 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=26640 $Y=20700 $dt=1
M40 97 A3 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=26660 $Y=4060 $dt=1
M41 VDD B3 96 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=27050 $Y=20700 $dt=1
M42 VDD B2 97 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=27070 $Y=4060 $dt=1
M43 24 96 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=27460 $Y=20700 $dt=1
M44 28 97 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=27480 $Y=4060 $dt=1
M45 98 A3 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=39760 $Y=20750 $dt=1
M46 VDD B3 98 VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=40170 $Y=20750 $dt=1
M47 31 98 VDD VDD g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=40580 $Y=20750 $dt=1
.ends mult
