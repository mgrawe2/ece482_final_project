************************************************************************
* auCdl Netlist:
* 
* Library Name:  ece482_final_project
* Top Cell Name: xor
* View Name:     schematic
* Netlisted on:  Nov 29 12:39:43 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: ece482_final_project
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv IN OUT VDD VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
MPM0 OUT IN VDD VDD g45p1svt m=1 l=45n w=240n
MNM0 OUT IN VSS VSS g45n1svt m=1 l=45n w=120n
.ENDS

************************************************************************
* Library Name: ece482_final_project
* Cell Name:    xor
* View Name:    schematic
************************************************************************

.SUBCKT xor A B B_bar OUT VDD VSS
*.PININFO A:I B:I B_bar:O OUT:O VDD:B VSS:B
MNM1 OUT A B_bar VSS g45n1svt m=1 l=45n w=120n
MNM0 A B_bar OUT VSS g45n1svt m=1 l=45n w=120n
MPM2 OUT A B VDD g45p1svt m=1 l=45n w=240n
MPM0 A B OUT VDD g45p1svt m=1 l=45n w=240n
XI0 B B_bar VDD VSS / inv
.ENDS

