* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : xor                                          *
* Netlisted  : Sat Nov 29 12:39:47 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764441582630                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764441582630 S_source_0 D_drain_1 3
** N=3 EP=3 FDC=1
M0 D_drain_1 3 S_source_0 S_source_0 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3034 scb=0.0125586 scc=0.000527096 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764441582630

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764441582631                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764441582631 S_source_0 D_drain_1 3 B
** N=5 EP=4 FDC=1
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=39.9325 scb=0.0377946 scc=0.00385132 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764441582631

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv IN OUT VDD VSS
** N=4 EP=4 FDC=2
X0 VSS OUT IN nmos1v_CDNS_764441582630 $T=-50 -540 0 0 $X=-470 $Y=-740
X1 VDD OUT IN VDD pmos1v_CDNS_764441582631 $T=-50 460 0 0 $X=-470 $Y=260
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764441582632                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764441582632 S_source_0 D_drain_1 S_source_2 B
** N=5 EP=4 FDC=2
M0 D_drain_1 S_source_2 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=48.7608 scb=0.0470044 scc=0.00589085 $X=0 $Y=0 $dt=1
M1 S_source_2 S_source_0 D_drain_1 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=56.1562 scb=0.0589139 scc=0.00666125 $X=410 $Y=0 $dt=1
.ends pmos1v_CDNS_764441582632

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764441582633                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764441582633 S_source_0 D_drain_1 S_source_2 4
** N=4 EP=4 FDC=2
M0 D_drain_1 S_source_2 S_source_0 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=5.12155 scb=0.00103813 scc=1.48881e-06 $X=0 $Y=0 $dt=0
M1 S_source_2 S_source_0 D_drain_1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=5.12155 scb=0.00103813 scc=1.48881e-06 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764441582633

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor A B B_Bar OUT VDD VSS
** N=6 EP=6 FDC=6
X5 B B_Bar VDD VSS inv $T=-790 -50 0 0 $X=-1590 $Y=-1230
X6 A OUT B VDD pmos1v_CDNS_764441582632 $T=660 1350 0 0 $X=240 $Y=1150
X7 A OUT B_Bar VSS nmos1v_CDNS_764441582633 $T=660 -340 0 0 $X=240 $Y=-540
.ends xor
