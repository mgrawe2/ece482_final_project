* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mult                                         *
* Netlisted  : Sun Nov 30 19:17:02 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764551816960                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764551816960 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764551816960

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764551816961                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764551816961 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764551816961

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764551816962                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764551816962 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764551816962

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764551816963                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764551816963 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_764551816963

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_764551816964                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_764551816964 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_764551816964

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764551816965                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764551816965 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764551816965

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764551816967                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764551816967 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764551816967

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764551816968                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764551816968 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764551816968

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764551816969                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764551816969 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764551816969

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7645518169610                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7645518169610 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7645518169610

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7645518169611                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7645518169611 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7645518169611

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7645518169612                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7645518169612 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7645518169612

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7645518169613                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7645518169613 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7645518169613

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7645518169614                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7645518169614 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7645518169614

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_7645518169615                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_7645518169615 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_7645518169615

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_7645518169616                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_7645518169616 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_7645518169616

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_7645518169617                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_7645518169617 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_7645518169617

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_7645518169618                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_7645518169618 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_7645518169618

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764551816960                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764551816960 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 3 1 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=7.55e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=0 $Y=0 $dt=1
M1 4 6 2 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=5.5e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=410 $Y=0 $dt=1
M2 5 7 4 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=3.45e-07 sca=30.7814 scb=0.0252726 scc=0.00362484 $X=820 $Y=0 $dt=1
M3 8 9 5 11 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=7.55e-07 sb=1.4e-07 sca=30.82 scb=0.02528 scc=0.00362484 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_764551816960

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764551816961                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764551816961 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_764551816961

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764551816962                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764551816962 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_764551816962

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764551816963                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764551816963 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764551816963

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
X0 4 3 1 nmos1v_CDNS_764551816962 $T=-50 -540 0 0 $X=-470 $Y=-740
X1 2 3 1 4 2 pmos1v_CDNS_764551816963 $T=-50 460 0 0 $X=-470 $Y=260
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764551816964                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764551816964 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764551816964

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764551816965                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764551816965 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=0 $Y=0 $dt=0
M1 3 1 2 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764551816965

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 5 M1_PO_CDNS_764551816960 $T=850 -1090 0 0 $X=750 $Y=-1450
X1 1 M1_PO_CDNS_764551816960 $T=850 2390 0 0 $X=750 $Y=2030
X2 4 M1_PO_CDNS_764551816960 $T=1260 650 0 0 $X=1160 $Y=290
X3 4 M2_M1_CDNS_764551816968 $T=360 650 0 0 $X=280 $Y=240
X4 4 M2_M1_CDNS_764551816968 $T=1260 650 0 0 $X=1180 $Y=240
X5 1 2 5 3 inv $T=-790 -50 0 0 $X=-1590 $Y=-1230
X6 4 6 1 3 2 pmos1v_CDNS_764551816964 $T=660 1350 0 0 $X=240 $Y=1150
X7 4 6 5 3 nmos1v_CDNS_764551816965 $T=660 -340 0 0 $X=240 $Y=-540
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 1 2 3 4 5 6 7 8 9 10
+ 13 14 15
** N=15 EP=13 FDC=22
X0 2 M1_PO_CDNS_764551816960 $T=790 -2720 0 0 $X=690 $Y=-3080
X1 8 M1_PO_CDNS_764551816960 $T=1490 -1360 0 0 $X=1390 $Y=-1720
X2 9 M1_PO_CDNS_764551816960 $T=1490 -160 0 0 $X=1390 $Y=-520
X3 9 M1_PO_CDNS_764551816960 $T=1900 -1360 0 0 $X=1800 $Y=-1720
X4 8 M1_PO_CDNS_764551816960 $T=1900 -160 0 0 $X=1800 $Y=-520
X5 5 M1_PO_CDNS_764551816960 $T=2310 -2720 0 0 $X=2210 $Y=-3080
X6 8 M2_M1_CDNS_764551816961 $T=-4410 -500 0 0 $X=-4490 $Y=-770
X7 6 M2_M1_CDNS_764551816961 $T=-610 -540 0 0 $X=-690 $Y=-810
X8 9 M2_M1_CDNS_764551816961 $T=-540 -2000 0 0 $X=-620 $Y=-2270
X9 10 M2_M1_CDNS_764551816961 $T=590 -90 0 0 $X=510 $Y=-360
X10 2 M2_M1_CDNS_764551816961 $T=790 -2710 0 0 $X=710 $Y=-2980
X11 8 M2_M1_CDNS_764551816961 $T=1490 -1390 0 0 $X=1410 $Y=-1660
X12 9 M2_M1_CDNS_764551816961 $T=1900 -1360 0 0 $X=1820 $Y=-1630
X13 8 M2_M1_CDNS_764551816961 $T=1900 -160 0 0 $X=1820 $Y=-430
X14 5 M2_M1_CDNS_764551816961 $T=2320 -2720 0 0 $X=2240 $Y=-2990
X15 10 M2_M1_CDNS_764551816961 $T=2510 -70 0 0 $X=2430 $Y=-340
X16 8 M3_M2_CDNS_764551816962 $T=-4410 -500 0 0 $X=-4490 $Y=-770
X17 6 M3_M2_CDNS_764551816962 $T=-610 -540 0 0 $X=-690 $Y=-810
X18 9 M3_M2_CDNS_764551816962 $T=-540 -2000 0 0 $X=-620 $Y=-2270
X19 10 M3_M2_CDNS_764551816962 $T=590 -90 0 0 $X=510 $Y=-360
X20 2 M3_M2_CDNS_764551816962 $T=790 -2710 0 0 $X=710 $Y=-2980
X21 9 M3_M2_CDNS_764551816962 $T=1900 -1360 0 0 $X=1820 $Y=-1630
X22 10 M3_M2_CDNS_764551816962 $T=2510 -70 0 0 $X=2430 $Y=-340
X23 3 M1_NWELL_CDNS_764551816963 $T=1520 1390 0 0 $X=1100 $Y=1090
X24 4 M1_PSUB_CDNS_764551816964 $T=1540 -3300 0 0 $X=1160 $Y=-3440
X25 3 M2_M1_CDNS_764551816965 $T=-6190 480 0 0 $X=-6410 $Y=350
X26 8 M2_M1_CDNS_764551816965 $T=-2450 -890 0 0 $X=-2670 $Y=-1020
X27 3 M2_M1_CDNS_764551816965 $T=-2390 480 0 0 $X=-2610 $Y=350
X28 3 M2_M1_CDNS_764551816965 $T=1530 1390 0 0 $X=1310 $Y=1260
X29 1 M3_M2_CDNS_764551816967 $T=-6990 -3990 0 0 $X=-7070 $Y=-4400
X30 5 M3_M2_CDNS_764551816967 $T=-4300 -3990 0 0 $X=-4380 $Y=-4400
X31 2 M3_M2_CDNS_764551816967 $T=-1030 -260 0 0 $X=-1110 $Y=-670
X32 6 M3_M2_CDNS_764551816967 $T=-600 2400 0 0 $X=-680 $Y=1990
X33 1 M2_M1_CDNS_764551816968 $T=-6990 -3990 0 0 $X=-7070 $Y=-4400
X34 5 M2_M1_CDNS_764551816968 $T=-4300 -3990 0 0 $X=-4380 $Y=-4400
X35 6 M2_M1_CDNS_764551816968 $T=-600 2400 0 0 $X=-680 $Y=1990
X36 2 M3_M2_CDNS_764551816969 $T=-7660 -2700 0 0 $X=-8020 $Y=-2830
X37 4 M3_M2_CDNS_764551816969 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X38 3 M3_M2_CDNS_764551816969 $T=3220 2330 0 0 $X=2860 $Y=2200
X39 7 M3_M2_CDNS_764551816969 $T=4650 0 0 0 $X=4290 $Y=-130
X40 2 M2_M1_CDNS_7645518169610 $T=-7660 -2700 0 0 $X=-8020 $Y=-2830
X41 4 M2_M1_CDNS_7645518169610 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X42 3 M2_M1_CDNS_7645518169610 $T=3220 2330 0 0 $X=2860 $Y=2200
X43 7 M2_M1_CDNS_7645518169610 $T=4650 0 0 0 $X=4290 $Y=-130
X44 4 M4_M3_CDNS_7645518169611 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X45 3 M4_M3_CDNS_7645518169611 $T=3220 2330 0 0 $X=2860 $Y=2200
X46 4 M5_M4_CDNS_7645518169612 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X47 3 M5_M4_CDNS_7645518169612 $T=3220 2330 0 0 $X=2860 $Y=2200
X48 4 M6_M5_CDNS_7645518169613 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X49 3 M6_M5_CDNS_7645518169613 $T=3220 2330 0 0 $X=2860 $Y=2200
X50 4 M7_M6_CDNS_7645518169614 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X51 3 M7_M6_CDNS_7645518169614 $T=3220 2330 0 0 $X=2860 $Y=2200
X52 4 M8_M7_CDNS_7645518169615 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X53 3 M8_M7_CDNS_7645518169615 $T=3220 2330 0 0 $X=2860 $Y=2200
X54 4 M9_M8_CDNS_7645518169616 $T=1570 -4010 0 0 $X=1210 $Y=-4140
X55 3 M9_M8_CDNS_7645518169616 $T=3220 2330 0 0 $X=2860 $Y=2200
X56 4 M10_M9_CDNS_7645518169617 $T=1590 -4010 0 0 $X=630 $Y=-4290
X57 3 M10_M9_CDNS_7645518169617 $T=3240 2340 0 0 $X=2280 $Y=2060
X58 4 M11_M10_CDNS_7645518169618 $T=1590 -4010 0 0 $X=630 $Y=-4290
X59 3 M11_M10_CDNS_7645518169618 $T=3240 2340 0 0 $X=2280 $Y=2060
X60 10 11 2 3 12 9 8 10 5 4
+ 3 pmos1v_CDNS_764551816960 $T=890 400 0 0 $X=470 $Y=200
X61 10 13 2 4 14 8 9 10 5 nmos1v_CDNS_764551816961 $T=890 -2160 0 0 $X=470 $Y=-2360
X62 10 3 7 4 inv $T=3440 20 0 0 $X=2640 $Y=-1160
X63 1 3 4 5 15 8 xor $T=-5190 -910 0 0 $X=-7060 $Y=-2360
X64 8 3 4 2 9 6 xor $T=-1390 -910 0 0 $X=-3260 $Y=-2360
M0 15 1 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.6083 scb=0.0129915 scc=0.000573075 $X=-6030 $Y=-1500 $dt=0
M1 9 8 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.6083 scb=0.0129915 scc=0.000573075 $X=-2230 $Y=-1500 $dt=0
M2 7 10 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=15.2291 scb=0.0163495 scc=0.00102074 $X=3390 $Y=-520 $dt=0
M3 15 1 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=38.1374 scb=0.0367153 scc=0.003591 $X=-6030 $Y=-500 $dt=1
M4 8 1 5 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-4530 $Y=440 $dt=1
M5 1 5 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-4120 $Y=440 $dt=1
M6 9 8 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=37.8604 scb=0.0362251 scc=0.00357304 $X=-2230 $Y=-500 $dt=1
M7 6 8 2 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-730 $Y=440 $dt=1
M8 8 2 6 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=43.4939 scb=0.0426265 scc=0.00546355 $X=-320 $Y=440 $dt=1
M9 7 10 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=28.8254 scb=0.0308995 scc=0.00229409 $X=3390 $Y=480 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_7645518169622                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_7645518169622 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_7645518169622

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764551816966                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764551816966 1 2 3 4 5 6 7 8
*.DEVICECLIMB
** N=8 EP=8 FDC=0
.ends pmos1v_CDNS_764551816966

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764551816967                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764551816967 1 2 3 4 5 6
** N=6 EP=6 FDC=3
M0 2 3 1 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 5 4 2 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 6 1 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
.ends nmos1v_CDNS_764551816967

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=3
X0 4 M1_PO_CDNS_764551816960 $T=-560 200 0 0 $X=-660 $Y=-160
X1 3 M1_PO_CDNS_764551816960 $T=-150 -970 0 0 $X=-250 $Y=-1330
X2 6 M1_PO_CDNS_764551816960 $T=260 -270 0 0 $X=160 $Y=-630
X3 4 M2_M1_CDNS_764551816961 $T=-560 200 0 0 $X=-640 $Y=-70
X4 3 M2_M1_CDNS_764551816961 $T=-150 -970 0 0 $X=-230 $Y=-1240
X5 4 M3_M2_CDNS_764551816962 $T=-560 200 0 0 $X=-640 $Y=-70
X6 3 M3_M2_CDNS_764551816962 $T=-150 -970 0 0 $X=-230 $Y=-1240
X7 1 M1_NWELL_CDNS_764551816963 $T=-10 1800 0 0 $X=-430 $Y=1500
X8 2 M1_PSUB_CDNS_764551816964 $T=-10 -2390 0 0 $X=-390 $Y=-2530
X9 3 M3_M2_CDNS_764551816967 $T=-1500 -4280 0 0 $X=-1580 $Y=-4690
X10 4 M3_M2_CDNS_764551816967 $T=-990 -4280 0 0 $X=-1070 $Y=-4690
X11 5 M3_M2_CDNS_764551816967 $T=990 2710 0 0 $X=910 $Y=2300
X12 3 M2_M1_CDNS_764551816968 $T=-1500 -4280 0 0 $X=-1580 $Y=-4690
X13 4 M2_M1_CDNS_764551816968 $T=-990 -4280 0 0 $X=-1070 $Y=-4690
X14 5 M2_M1_CDNS_764551816968 $T=990 2710 0 0 $X=910 $Y=2300
X15 1 M3_M2_CDNS_764551816969 $T=-640 2480 0 0 $X=-1000 $Y=2350
X16 2 M3_M2_CDNS_764551816969 $T=680 -3080 0 0 $X=320 $Y=-3210
X17 1 M2_M1_CDNS_7645518169610 $T=-640 2480 0 0 $X=-1000 $Y=2350
X18 2 M2_M1_CDNS_7645518169610 $T=680 -3080 0 0 $X=320 $Y=-3210
X19 1 M4_M3_CDNS_7645518169611 $T=-640 2480 0 0 $X=-1000 $Y=2350
X20 2 M4_M3_CDNS_7645518169611 $T=680 -3080 0 0 $X=320 $Y=-3210
X21 1 M5_M4_CDNS_7645518169612 $T=-640 2480 0 0 $X=-1000 $Y=2350
X22 2 M5_M4_CDNS_7645518169612 $T=680 -3080 0 0 $X=320 $Y=-3210
X23 1 M6_M5_CDNS_7645518169613 $T=-640 2480 0 0 $X=-1000 $Y=2350
X24 2 M6_M5_CDNS_7645518169613 $T=680 -3080 0 0 $X=320 $Y=-3210
X25 1 M7_M6_CDNS_7645518169614 $T=-640 2480 0 0 $X=-1000 $Y=2350
X26 2 M7_M6_CDNS_7645518169614 $T=680 -3080 0 0 $X=320 $Y=-3210
X27 1 M8_M7_CDNS_7645518169615 $T=-640 2480 0 0 $X=-1000 $Y=2350
X28 2 M8_M7_CDNS_7645518169615 $T=680 -3080 0 0 $X=320 $Y=-3210
X29 1 M9_M8_CDNS_7645518169616 $T=-640 2480 0 0 $X=-1000 $Y=2350
X30 2 M9_M8_CDNS_7645518169616 $T=680 -3080 0 0 $X=320 $Y=-3210
X31 1 M10_M9_CDNS_7645518169617 $T=-630 2470 0 0 $X=-1590 $Y=2190
X32 2 M10_M9_CDNS_7645518169617 $T=700 -3080 0 0 $X=-260 $Y=-3360
X33 1 M11_M10_CDNS_7645518169622 $T=-630 2470 0 0 $X=-1590 $Y=2190
X34 2 M11_M10_CDNS_7645518169622 $T=700 -3080 0 0 $X=-260 $Y=-3360
X35 1 6 4 3 1 5 2 1 pmos1v_CDNS_764551816966 $T=-460 820 0 0 $X=-880 $Y=620
X36 6 7 4 3 2 5 nmos1v_CDNS_764551816967 $T=-460 -1890 0 0 $X=-880 $Y=-2090
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 7
** N=9 EP=7 FDC=12
X0 5 M2_M1_CDNS_764551816961 $T=-1450 460 0 0 $X=-1530 $Y=190
X1 5 M3_M2_CDNS_764551816962 $T=-1450 460 0 0 $X=-1530 $Y=190
X2 1 M3_M2_CDNS_764551816967 $T=-4170 -2510 0 0 $X=-4250 $Y=-2920
X3 4 M3_M2_CDNS_764551816967 $T=-1860 -2510 0 0 $X=-1940 $Y=-2920
X4 4 M3_M2_CDNS_764551816967 $T=-1860 720 0 0 $X=-1940 $Y=310
X5 5 M3_M2_CDNS_764551816967 $T=-1450 3410 0 0 $X=-1530 $Y=3000
X6 1 M2_M1_CDNS_764551816968 $T=-4170 -2510 0 0 $X=-4250 $Y=-2920
X7 1 M2_M1_CDNS_764551816968 $T=-4170 440 0 0 $X=-4250 $Y=30
X8 4 M2_M1_CDNS_764551816968 $T=-1860 -2510 0 0 $X=-1940 $Y=-2920
X9 5 M2_M1_CDNS_764551816968 $T=-1450 3410 0 0 $X=-1530 $Y=3000
X10 2 M2_M1_CDNS_7645518169610 $T=-3220 1460 0 0 $X=-3580 $Y=1330
X11 2 M2_M1_CDNS_7645518169610 $T=620 2430 0 0 $X=260 $Y=2300
X12 1 2 3 4 7 5 xor $T=-2220 70 0 0 $X=-4090 $Y=-1380
X13 2 3 1 4 6 8 9 and2 $T=630 630 0 0 $X=-960 $Y=-4060
M0 7 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.9282 scb=0.0134361 scc=0.000622896 $X=-3060 $Y=-520 $dt=0
M1 7 1 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=36.6317 scb=0.035909 scc=0.00335548 $X=-3060 $Y=480 $dt=1
M2 5 1 4 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=-1560 $Y=1420 $dt=1
M3 1 4 5 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=-1150 $Y=1420 $dt=1
M4 8 4 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=26.2992 scb=0.0240146 scc=0.00255754 $X=170 $Y=1450 $dt=1
M5 2 1 8 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=28.7383 scb=0.0277231 scc=0.00260208 $X=580 $Y=1450 $dt=1
M6 6 8 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=39.2498 scb=0.0428135 scc=0.00408073 $X=990 $Y=1450 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mult                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mult 35 37 41 44 34 39 42 45 36 48
+ 49 50 19 26 32 33 3 4
** N=142 EP=18 FDC=320
X0 1 2 3 4 5 6 7 52 53 54
+ 107 108 51 full_adder $T=-5100 -5060 0 0 $X=-13120 $Y=-9460
X1 8 9 3 4 10 11 12 56 57 58
+ 109 110 55 full_adder $T=7620 11130 0 0 $X=-400 $Y=6730
X2 13 7 3 4 14 10 15 60 61 62
+ 111 112 59 full_adder $T=8320 -5030 0 0 $X=300 $Y=-9430
X3 16 17 3 4 18 19 20 64 65 66
+ 113 114 63 full_adder $T=20720 27820 0 0 $X=12700 $Y=23420
X4 21 12 3 4 22 18 23 68 69 70
+ 115 116 67 full_adder $T=21270 11120 0 0 $X=13250 $Y=6720
X5 24 20 3 4 25 26 27 72 73 74
+ 117 118 71 full_adder $T=34370 27810 0 0 $X=26350 $Y=23410
X6 28 23 3 4 29 25 30 76 77 78
+ 119 120 75 full_adder $T=35050 11120 0 0 $X=27030 $Y=6720
X7 31 27 3 4 30 32 33 80 81 82
+ 121 122 79 full_adder $T=48150 27810 0 0 $X=40130 $Y=23410
X8 3 4 34 35 36 83 123 and2 $T=-26670 -21260 0 0 $X=-28260 $Y=-25950
X9 3 4 34 37 38 84 124 and2 $T=-22280 -21130 0 0 $X=-23870 $Y=-25820
X10 3 4 39 35 40 85 125 and2 $T=-18840 -12210 0 0 $X=-20430 $Y=-16900
X11 3 4 34 41 5 86 126 and2 $T=-13020 -21220 0 0 $X=-14610 $Y=-25910
X12 3 4 42 35 43 87 127 and2 $T=-12210 3290 0 0 $X=-13800 $Y=-1400
X13 3 4 39 37 1 88 128 and2 $T=-10040 -12640 0 0 $X=-11630 $Y=-17330
X14 3 4 42 37 8 89 129 and2 $T=400 3630 0 0 $X=-1190 $Y=-1060
X15 3 4 34 44 14 90 130 and2 $T=540 -21460 0 0 $X=-1050 $Y=-26150
X16 3 4 45 35 46 91 131 and2 $T=890 19980 0 0 $X=-700 $Y=15290
X17 3 4 39 41 13 92 132 and2 $T=3520 -12410 0 0 $X=1930 $Y=-17100
X18 3 4 45 37 16 93 133 and2 $T=13500 20320 0 0 $X=11910 $Y=15630
X19 3 4 42 41 21 94 134 and2 $T=14000 3190 0 0 $X=12410 $Y=-1500
X20 3 4 39 44 47 95 135 and2 $T=15640 -12550 0 0 $X=14050 $Y=-17240
X21 3 4 45 41 24 96 136 and2 $T=27100 19880 0 0 $X=25510 $Y=15190
X22 3 4 42 44 28 97 137 and2 $T=27120 3240 0 0 $X=25530 $Y=-1450
X23 3 4 45 44 31 98 138 and2 $T=40220 19930 0 0 $X=38630 $Y=15240
X24 40 3 4 38 48 2 99 half_adder $T=-15990 -5900 0 0 $X=-20240 $Y=-9960
X25 43 3 4 6 49 9 101 half_adder $T=-7050 9650 0 0 $X=-11300 $Y=5590
X26 46 3 4 11 50 17 103 half_adder $T=6050 26340 0 0 $X=1800 $Y=22280
X27 15 3 4 47 22 29 105 half_adder $T=18470 -5780 0 0 $X=14220 $Y=-9840
M0 83 35 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-27130 $Y=-20440 $dt=1
M1 3 34 83 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-26720 $Y=-20440 $dt=1
M2 36 83 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-26310 $Y=-20440 $dt=1
M3 84 37 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-22740 $Y=-20310 $dt=1
M4 3 34 84 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-22330 $Y=-20310 $dt=1
M5 38 84 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-21920 $Y=-20310 $dt=1
M6 85 35 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-19300 $Y=-11390 $dt=1
M7 3 39 85 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-18890 $Y=-11390 $dt=1
M8 40 85 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-18480 $Y=-11390 $dt=1
M9 86 41 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-13480 $Y=-20400 $dt=1
M10 3 34 86 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-13070 $Y=-20400 $dt=1
M11 87 35 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-12670 $Y=4110 $dt=1
M12 5 86 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-12660 $Y=-20400 $dt=1
M13 3 42 87 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-12260 $Y=4110 $dt=1
M14 43 87 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-11850 $Y=4110 $dt=1
M15 88 37 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-10500 $Y=-11820 $dt=1
M16 3 39 88 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=-10090 $Y=-11820 $dt=1
M17 1 88 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=-9680 $Y=-11820 $dt=1
M18 89 37 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=-60 $Y=4450 $dt=1
M19 90 44 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=80 $Y=-20640 $dt=1
M20 3 42 89 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=350 $Y=4450 $dt=1
M21 91 35 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=430 $Y=20800 $dt=1
M22 3 34 90 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=490 $Y=-20640 $dt=1
M23 8 89 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=760 $Y=4450 $dt=1
M24 3 45 91 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=840 $Y=20800 $dt=1
M25 14 90 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=900 $Y=-20640 $dt=1
M26 46 91 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=1250 $Y=20800 $dt=1
M27 92 41 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=3060 $Y=-11590 $dt=1
M28 3 39 92 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=3470 $Y=-11590 $dt=1
M29 13 92 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=3880 $Y=-11590 $dt=1
M30 93 37 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=13040 $Y=21140 $dt=1
M31 3 45 93 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=13450 $Y=21140 $dt=1
M32 94 41 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=13540 $Y=4010 $dt=1
M33 16 93 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=13860 $Y=21140 $dt=1
M34 3 42 94 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=13950 $Y=4010 $dt=1
M35 21 94 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=14360 $Y=4010 $dt=1
M36 95 44 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=15180 $Y=-11730 $dt=1
M37 3 39 95 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=15590 $Y=-11730 $dt=1
M38 47 95 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=16000 $Y=-11730 $dt=1
M39 96 41 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=26640 $Y=20700 $dt=1
M40 97 44 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=26660 $Y=4060 $dt=1
M41 3 45 96 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=27050 $Y=20700 $dt=1
M42 3 42 97 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=27070 $Y=4060 $dt=1
M43 24 96 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=27460 $Y=20700 $dt=1
M44 28 97 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=27480 $Y=4060 $dt=1
M45 98 44 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=39760 $Y=20750 $dt=1
M46 3 45 98 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=40170 $Y=20750 $dt=1
M47 31 98 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=40580 $Y=20750 $dt=1
.ends mult
