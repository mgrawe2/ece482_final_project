* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : half_adder                                   *
* Netlisted  : Sun Nov 30 14:03:59 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764533033910                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764533033910 S_source_0 D_drain_1 3
** N=3 EP=3 FDC=1
M0 D_drain_1 3 S_source_0 S_source_0 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.9282 scb=0.0134361 scc=0.000622896 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764533033910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764533033911                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764533033911 S_source_0 D_drain_1 3 B
** N=5 EP=4 FDC=1
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=36.6317 scb=0.035909 scc=0.00335548 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764533033911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv VDD IN OUT VSS
** N=4 EP=4 FDC=2
X0 VSS OUT IN nmos1v_CDNS_764533033910 $T=-50 -540 0 0 $X=-470 $Y=-740
X1 VDD OUT IN VDD pmos1v_CDNS_764533033911 $T=-50 460 0 0 $X=-470 $Y=260
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764533033912                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764533033912 S_source_0 D_drain_1 S_source_2 B
** N=5 EP=4 FDC=2
M0 D_drain_1 S_source_2 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=0 $Y=0 $dt=1
M1 S_source_2 S_source_0 D_drain_1 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=410 $Y=0 $dt=1
.ends pmos1v_CDNS_764533033912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764533033913                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764533033913 S_source_0 D_drain_1 S_source_2 4
** N=4 EP=4 FDC=2
M0 D_drain_1 S_source_2 S_source_0 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=0 $Y=0 $dt=0
M1 S_source_2 S_source_0 D_drain_1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764533033913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor VDD VSS B B_Bar 5 OUT
** N=6 EP=6 FDC=6
X5 VDD B B_Bar VSS inv $T=-790 -50 0 0 $X=-1590 $Y=-1230
X6 5 OUT B VDD pmos1v_CDNS_764533033912 $T=660 1350 0 0 $X=240 $Y=1150
X7 5 OUT B_Bar VSS nmos1v_CDNS_764533033913 $T=660 -340 0 0 $X=240 $Y=-540
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764533033914                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764533033914 S_source_0 D_drain_1 3 4 S_source_2 D_drain_3 B
** N=8 EP=7 FDC=3
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=26.2992 scb=0.0240146 scc=0.00255754 $X=0 $Y=0 $dt=1
M1 S_source_2 4 D_drain_1 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=28.7383 scb=0.0277231 scc=0.00260208 $X=410 $Y=0 $dt=1
M2 D_drain_3 D_drain_1 S_source_2 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=39.2498 scb=0.0428135 scc=0.00408073 $X=820 $Y=0 $dt=1
.ends pmos1v_CDNS_764533033914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764533033915                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764533033915 S_source_0 D_drain_1 3 4 S_source_2 D_drain_3
** N=6 EP=6 FDC=3
M0 D_drain_1 3 S_source_0 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 S_source_2 4 D_drain_1 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 D_drain_3 S_source_0 S_source_2 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
.ends nmos1v_CDNS_764533033915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 VDD VSS A B OUT
** N=7 EP=5 FDC=6
X33 VDD 6 A B VDD OUT VDD pmos1v_CDNS_764533033914 $T=-460 820 0 0 $X=-880 $Y=620
X34 6 7 A B VSS OUT nmos1v_CDNS_764533033915 $T=-460 -1890 0 0 $X=-880 $Y=-2090
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder A B Co S VDD VSS
** N=9 EP=6 FDC=12
X12 VDD VSS B 6 A S xor $T=-2220 70 0 0 $X=-4090 $Y=-1380
X13 VDD VSS A B Co and2 $T=630 630 0 0 $X=-960 $Y=-4060
.ends half_adder
