* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : and2                                         *
* Netlisted  : Sun Nov 30 13:51:59 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764532313970                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764532313970 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764532313970

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764532313973                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764532313973 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764532313973

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764532313974                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764532313974 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764532313974

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_764532313975                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_764532313975 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_764532313975

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_764532313976                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_764532313976 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_764532313976

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_764532313977                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_764532313977 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_764532313977

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_764532313978                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_764532313978 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_764532313978

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_764532313979                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_764532313979 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_764532313979

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_7645323139710                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_7645323139710 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_7645323139710

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_7645323139711                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_7645323139711 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_7645323139711

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_7645323139712                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_7645323139712 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_7645323139712

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7645323139713                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7645323139713 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7645323139713

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7645323139714                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7645323139714 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7645323139714

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7645323139715                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7645323139715 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7645323139715

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764532313970                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764532313970 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=3
M0 2 3 1 8 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=0 $Y=0 $dt=1
M1 5 4 2 8 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=410 $Y=0 $dt=1
M2 6 2 5 8 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=820 $Y=0 $dt=1
.ends pmos1v_CDNS_764532313970

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764532313971                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764532313971 1 2 3 4 5 6
** N=6 EP=6 FDC=3
M0 2 3 1 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 5 4 2 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 6 1 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
.ends nmos1v_CDNS_764532313971

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 6 4 5
** N=7 EP=5 FDC=6
X0 1 M1_PO_CDNS_764532313970 $T=-560 200 0 0 $X=-660 $Y=-160
X1 2 M1_PO_CDNS_764532313970 $T=-150 -970 0 0 $X=-250 $Y=-1330
X2 3 M1_PO_CDNS_764532313970 $T=260 -270 0 0 $X=160 $Y=-630
X3 4 M3_M2_CDNS_764532313973 $T=-650 2430 0 0 $X=-1010 $Y=2300
X4 5 M3_M2_CDNS_764532313973 $T=680 -3080 0 0 $X=320 $Y=-3210
X5 4 M2_M1_CDNS_764532313974 $T=-650 2430 0 0 $X=-1010 $Y=2300
X6 5 M2_M1_CDNS_764532313974 $T=680 -3080 0 0 $X=320 $Y=-3210
X7 4 M4_M3_CDNS_764532313975 $T=-650 2430 0 0 $X=-1010 $Y=2300
X8 5 M4_M3_CDNS_764532313975 $T=680 -3080 0 0 $X=320 $Y=-3210
X9 4 M5_M4_CDNS_764532313976 $T=-650 2430 0 0 $X=-1010 $Y=2300
X10 5 M5_M4_CDNS_764532313976 $T=680 -3080 0 0 $X=320 $Y=-3210
X11 4 M6_M5_CDNS_764532313977 $T=-650 2430 0 0 $X=-1010 $Y=2300
X12 5 M6_M5_CDNS_764532313977 $T=680 -3080 0 0 $X=320 $Y=-3210
X13 4 M7_M6_CDNS_764532313978 $T=-650 2430 0 0 $X=-1010 $Y=2300
X14 5 M7_M6_CDNS_764532313978 $T=680 -3080 0 0 $X=320 $Y=-3210
X15 4 M8_M7_CDNS_764532313979 $T=-650 2430 0 0 $X=-1010 $Y=2300
X16 5 M8_M7_CDNS_764532313979 $T=680 -3080 0 0 $X=320 $Y=-3210
X17 4 M9_M8_CDNS_7645323139710 $T=-650 2430 0 0 $X=-1010 $Y=2300
X18 5 M9_M8_CDNS_7645323139710 $T=680 -3080 0 0 $X=320 $Y=-3210
X19 4 M10_M9_CDNS_7645323139711 $T=-630 2430 0 0 $X=-1590 $Y=2150
X20 5 M10_M9_CDNS_7645323139711 $T=700 -3080 0 0 $X=-260 $Y=-3360
X21 4 M11_M10_CDNS_7645323139712 $T=-630 2430 0 0 $X=-1590 $Y=2150
X22 5 M11_M10_CDNS_7645323139712 $T=700 -3080 0 0 $X=-260 $Y=-3360
X23 2 M2_M1_CDNS_7645323139713 $T=-1500 -4280 0 0 $X=-1580 $Y=-4690
X24 1 M2_M1_CDNS_7645323139713 $T=-990 -4280 0 0 $X=-1070 $Y=-4690
X25 6 M2_M1_CDNS_7645323139713 $T=990 2710 0 0 $X=910 $Y=2300
X26 2 M3_M2_CDNS_7645323139714 $T=-1500 -4280 0 0 $X=-1580 $Y=-4690
X27 1 M3_M2_CDNS_7645323139714 $T=-990 -4280 0 0 $X=-1070 $Y=-4690
X28 6 M3_M2_CDNS_7645323139714 $T=990 2710 0 0 $X=910 $Y=2300
X29 1 M2_M1_CDNS_7645323139715 $T=-560 200 0 0 $X=-640 $Y=-70
X30 2 M2_M1_CDNS_7645323139715 $T=-150 -970 0 0 $X=-230 $Y=-1240
X31 4 3 1 2 4 6 5 4 pmos1v_CDNS_764532313970 $T=-460 820 0 0 $X=-880 $Y=620
X32 3 7 1 2 5 6 nmos1v_CDNS_764532313971 $T=-460 -1890 0 0 $X=-880 $Y=-2090
.ends and2
