* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pipeline_mult                                *
* Netlisted  : Sun Dec  7 19:50:41 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_765158635880                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_765158635880 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_765158635880

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765158635881                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765158635881 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765158635881

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765158635882                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765158635882 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765158635882

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765158635883                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765158635883 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765158635883

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765158635884                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765158635884 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765158635884

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765158635885                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765158635885 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765158635885

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765158635886                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765158635886 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765158635886

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765158635887                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765158635887 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765158635887

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765158635888                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765158635888 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765158635888

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765158635889                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765158635889 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765158635889

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_7651586358810                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_7651586358810 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_7651586358810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7651586358811                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7651586358811 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7651586358811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7651586358812                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7651586358812 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7651586358812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7651586358813                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7651586358813 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7651586358813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651586358814                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651586358814 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651586358814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651586358815                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651586358815 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651586358815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_7651586358816                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_7651586358816 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_7651586358816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651586358817                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651586358817 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651586358817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651586358818                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651586358818 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651586358818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7651586358819                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7651586358819 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7651586358819

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651586358820                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651586358820 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651586358820

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_7651586358821                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_7651586358821 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_7651586358821

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651586358822                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651586358822 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651586358822

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651586358823                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651586358823 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651586358823

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765158635880                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765158635880 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765158635880

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158635881                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158635881 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765158635881

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158635882                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158635882 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_765158635882

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: c2mos                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt c2mos 1 2 3 4 5 6 7 8 11 12
*.DEVICECLIMB
** N=12 EP=10 FDC=9
X0 1 M2_M1_CDNS_765158635885 $T=480 1970 0 90 $X=350 $Y=1890
X1 7 M2_M1_CDNS_765158635885 $T=1070 1420 0 90 $X=940 $Y=1340
X2 1 M2_M1_CDNS_765158635885 $T=3650 1970 0 90 $X=3520 $Y=1890
X3 7 M2_M1_CDNS_765158635885 $T=3660 1420 0 90 $X=3530 $Y=1340
X4 8 M2_M1_CDNS_765158635885 $T=4060 1720 0 90 $X=3930 $Y=1640
X5 8 M2_M1_CDNS_765158635885 $T=5220 1720 0 90 $X=5090 $Y=1640
X6 1 M2_M1_CDNS_765158635885 $T=5960 2040 0 90 $X=5830 $Y=1960
X7 7 M2_M1_CDNS_765158635885 $T=6620 1970 0 90 $X=6490 $Y=1890
X8 1 M1_PO_CDNS_7651586358822 $T=3660 1980 0 90 $X=3540 $Y=1880
X9 7 M1_PO_CDNS_7651586358822 $T=3670 1420 0 90 $X=3550 $Y=1320
X10 8 M1_PO_CDNS_7651586358822 $T=5210 1720 0 90 $X=5090 $Y=1620
X11 7 M1_PO_CDNS_7651586358822 $T=6630 1980 0 90 $X=6510 $Y=1880
X12 1 M1_PO_CDNS_7651586358822 $T=6660 1400 0 90 $X=6540 $Y=1300
X13 1 M1_PO_CDNS_7651586358823 $T=530 1970 0 0 $X=310 $Y=1850
X14 4 M1_PO_CDNS_7651586358823 $T=2110 1720 0 0 $X=1890 $Y=1600
X15 6 M1_PO_CDNS_7651586358823 $T=8090 1590 0 0 $X=7870 $Y=1470
X16 2 7 1 3 2 pmos1v_CDNS_765158635880 $T=750 2360 0 0 $X=330 $Y=2160
X17 2 9 4 3 2 pmos1v_CDNS_765158635880 $T=2240 2360 0 0 $X=1820 $Y=2160
X18 9 8 1 3 2 pmos1v_CDNS_765158635880 $T=3740 2350 0 0 $X=3320 $Y=2150
X19 2 10 8 3 2 pmos1v_CDNS_765158635880 $T=5230 2360 0 0 $X=4810 $Y=2160
X20 10 5 7 3 2 pmos1v_CDNS_765158635880 $T=6720 2340 0 0 $X=6300 $Y=2140
X21 3 1 7 3 nmos1v_CDNS_765158635881 $T=750 650 0 0 $X=330 $Y=450
X22 3 4 11 3 nmos1v_CDNS_765158635881 $T=2240 650 0 0 $X=1820 $Y=450
X23 11 7 8 3 nmos1v_CDNS_765158635881 $T=3750 650 0 0 $X=3330 $Y=450
X24 3 8 12 3 nmos1v_CDNS_765158635881 $T=5230 650 0 0 $X=4810 $Y=450
X25 12 1 5 3 nmos1v_CDNS_765158635881 $T=6720 650 0 0 $X=6300 $Y=450
X26 5 3 6 nmos1v_CDNS_765158635882 $T=8210 170 0 0 $X=7790 $Y=-30
M0 11 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=2240 $Y=650 $dt=0
M1 8 7 11 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=3750 $Y=650 $dt=0
M2 12 8 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=5230 $Y=650 $dt=0
M3 5 1 12 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=6720 $Y=650 $dt=0
M4 7 1 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.27 scb=0.0231774 scc=0.00199917 $X=750 $Y=2360 $dt=1
M5 9 4 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=2240 $Y=2360 $dt=1
M6 8 1 9 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.7063 scb=0.016025 scc=0.00198503 $X=3740 $Y=2350 $dt=1
M7 10 8 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=5230 $Y=2360 $dt=1
M8 5 7 10 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.6749 scb=0.0214174 scc=0.0021813 $X=6720 $Y=2340 $dt=1
.ends c2mos

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_7651586358828                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_7651586358828 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_7651586358828

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651586358829                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651586358829 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651586358829

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_7651586358830                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_7651586358830 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_7651586358830

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651586358831                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651586358831 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651586358831

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158635883                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158635883 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765158635883

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765158635884                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765158635884 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_765158635884

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158635885                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158635885 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765158635885

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X0 2 M1_NWELL_CDNS_7651586358828 $T=190 2570 0 0 $X=-230 $Y=2270
X1 4 M1_PSUB_CDNS_7651586358830 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 1 M1_PO_CDNS_7651586358831 $T=-160 30 0 0 $X=-260 $Y=-330
X3 2 3 1 2 4 2 pmos1v_CDNS_765158635884 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 3 1 4 4 nmos1v_CDNS_765158635885 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=9
X0 2 M1_NWELL_CDNS_7651586358828 $T=-1350 2870 0 0 $X=-1770 $Y=2570
X1 6 M2_M1_CDNS_7651586358829 $T=-2410 -1220 0 0 $X=-2490 $Y=-1470
X2 7 M2_M1_CDNS_7651586358829 $T=-2000 1650 0 0 $X=-2080 $Y=1400
X3 6 M2_M1_CDNS_7651586358829 $T=-1590 -1220 0 0 $X=-1670 $Y=-1470
X4 6 M2_M1_CDNS_7651586358829 $T=-1110 -1220 0 0 $X=-1190 $Y=-1470
X5 7 M2_M1_CDNS_7651586358829 $T=-700 1650 0 0 $X=-780 $Y=1400
X6 6 M2_M1_CDNS_7651586358829 $T=-290 -1220 0 0 $X=-370 $Y=-1470
X7 4 M1_PSUB_CDNS_7651586358830 $T=-700 -2440 0 0 $X=-1080 $Y=-2580
X8 1 M1_PO_CDNS_7651586358831 $T=-2350 360 0 0 $X=-2450 $Y=0
X9 3 M1_PO_CDNS_7651586358831 $T=-1050 60 0 0 $X=-1150 $Y=-300
X10 6 6 7 1 4 nmos1v_CDNS_765158635883 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 6 6 4 3 4 nmos1v_CDNS_765158635883 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X12 2 7 1 2 4 2 pmos1v_CDNS_765158635884 $T=-2250 930 0 0 $X=-2670 $Y=730
X13 2 7 3 2 4 2 pmos1v_CDNS_765158635884 $T=-950 930 0 0 $X=-1370 $Y=730
X14 7 2 5 4 inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 2 3 7 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M1 5 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M2 2 7 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651586358826                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651586358826 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651586358826

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651586358827                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651586358827 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651586358827

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X0 1 M1_PO_CDNS_7651586358822 $T=-450 10 0 0 $X=-550 $Y=-110
X1 1 M1_PO_CDNS_7651586358822 $T=-450 1890 0 0 $X=-550 $Y=1770
X2 4 M1_PO_CDNS_7651586358822 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X3 1 M1_PO_CDNS_7651586358822 $T=-40 1890 0 0 $X=-140 $Y=1770
X4 6 M1_PO_CDNS_7651586358822 $T=850 -980 0 0 $X=750 $Y=-1100
X5 4 M1_PO_CDNS_7651586358823 $T=-250 -840 0 0 $X=-470 $Y=-960
X6 6 M2_M1_CDNS_7651586358826 $T=-30 -450 0 0 $X=-160 $Y=-580
X7 5 M2_M1_CDNS_7651586358826 $T=1330 -190 0 0 $X=1200 $Y=-320
X8 6 M2_M1_CDNS_7651586358827 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X9 6 M2_M1_CDNS_7651586358827 $T=-250 380 0 0 $X=-380 $Y=250
X10 5 M2_M1_CDNS_7651586358829 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X11 5 M2_M1_CDNS_7651586358829 $T=-660 950 0 0 $X=-740 $Y=700
X12 5 M2_M1_CDNS_7651586358829 $T=160 -1560 0 0 $X=80 $Y=-1810
X13 5 M2_M1_CDNS_7651586358829 $T=160 950 0 0 $X=80 $Y=700
X14 5 M2_M1_CDNS_7651586358829 $T=1050 -1560 0 0 $X=970 $Y=-1810
X15 5 M2_M1_CDNS_7651586358829 $T=1050 950 0 0 $X=970 $Y=700
X16 5 6 1 5 3 2 pmos1v_CDNS_765158635884 $T=-500 230 0 0 $X=-920 $Y=30
X17 1 5 6 1 3 2 pmos1v_CDNS_765158635884 $T=800 230 0 0 $X=380 $Y=30
X18 5 6 4 5 3 nmos1v_CDNS_765158635885 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X19 4 5 6 4 3 nmos1v_CDNS_765158635885 $T=800 -1920 0 0 $X=380 $Y=-2120
X20 1 2 4 3 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
M0 5 1 6 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 5 6 1 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 1 6 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 7
** N=9 EP=7 FDC=24
X0 1 M3_M2_CDNS_765158635884 $T=2760 3570 0 0 $X=2680 $Y=3440
X1 2 M3_M2_CDNS_765158635884 $T=4630 3110 0 0 $X=4550 $Y=2980
X2 6 M3_M2_CDNS_765158635884 $T=9970 3310 0 0 $X=9890 $Y=3180
X3 5 M3_M2_CDNS_765158635884 $T=10180 2730 0 0 $X=10100 $Y=2600
X4 6 M2_M1_CDNS_765158635885 $T=9970 3310 0 0 $X=9890 $Y=3180
X5 5 M2_M1_CDNS_765158635885 $T=10180 2730 0 0 $X=10100 $Y=2600
X6 1 M2_M1_CDNS_7651586358826 $T=2760 2580 0 0 $X=2630 $Y=2450
X7 1 M2_M1_CDNS_7651586358826 $T=7960 2810 0 0 $X=7830 $Y=2680
X8 5 M2_M1_CDNS_7651586358827 $T=6360 3430 0 0 $X=6230 $Y=3300
X9 2 4 1 3 6 9 8 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X10 1 4 3 7 5 2 xor $T=4660 3560 0 0 $X=2440 $Y=1000
M0 7 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2860 $Y=3790 $dt=1
M1 4 1 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3270 $Y=3790 $dt=1
M2 2 1 5 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4160 $Y=3790 $dt=1
M3 8 2 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6760 $Y=3790 $dt=1
M4 4 2 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7170 $Y=3790 $dt=1
M5 8 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8060 $Y=3790 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651586358835                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651586358835 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651586358835

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158635886                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158635886 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_765158635886

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765158635887                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765158635887 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_765158635887

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=8
X0 1 M2_M1_CDNS_765158635885 $T=-830 -970 0 0 $X=-910 $Y=-1100
X1 2 M2_M1_CDNS_765158635885 $T=-220 -60 0 0 $X=-300 $Y=-190
X2 2 M2_M1_CDNS_765158635885 $T=200 730 0 0 $X=120 $Y=600
X3 1 M2_M1_CDNS_765158635885 $T=810 -970 0 0 $X=730 $Y=-1100
X4 2 M1_PO_CDNS_7651586358822 $T=-220 -60 0 0 $X=-320 $Y=-180
X5 5 M1_PO_CDNS_7651586358822 $T=-210 730 0 0 $X=-310 $Y=610
X6 5 M1_PO_CDNS_7651586358822 $T=190 -60 0 0 $X=90 $Y=-180
X7 2 M1_PO_CDNS_7651586358822 $T=200 730 0 0 $X=100 $Y=610
X8 4 M1_NWELL_CDNS_7651586358828 $T=-10 2990 0 0 $X=-430 $Y=2690
X9 6 M1_PSUB_CDNS_7651586358830 $T=0 -1600 0 0 $X=-380 $Y=-1740
X10 3 M1_PO_CDNS_7651586358831 $T=-590 550 0 0 $X=-690 $Y=190
X11 7 M1_PO_CDNS_7651586358831 $T=570 550 0 0 $X=470 $Y=190
X12 1 8 3 6 9 2 5 1 7 nmos1v_CDNS_765158635886 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 1 10 4 3 5 11 1 2 7 6
+ 4 pmos1v_CDNS_765158635887 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 1 2 3 4 5 6 7 8 9 10
+ 11
** N=15 EP=11 FDC=36
X0 2 M4_M3_CDNS_765158635882 $T=6980 3080 0 0 $X=6900 $Y=2950
X1 2 M4_M3_CDNS_765158635882 $T=10140 2970 0 0 $X=10060 $Y=2840
X2 1 M3_M2_CDNS_765158635884 $T=2270 3860 0 0 $X=2190 $Y=3730
X3 2 M3_M2_CDNS_765158635884 $T=5790 3080 0 0 $X=5710 $Y=2950
X4 6 M3_M2_CDNS_765158635884 $T=9120 4760 0 0 $X=9040 $Y=4630
X5 2 M3_M2_CDNS_765158635884 $T=11410 2940 0 0 $X=11330 $Y=2810
X6 7 M3_M2_CDNS_765158635884 $T=12920 3510 0 0 $X=12840 $Y=3380
X7 2 M2_M1_CDNS_765158635885 $T=5250 3070 0 0 $X=5170 $Y=2940
X8 8 M2_M1_CDNS_765158635885 $T=9530 2380 0 0 $X=9450 $Y=2250
X9 9 M2_M1_CDNS_765158635885 $T=9530 5090 0 0 $X=9450 $Y=4960
X10 4 M2_M1_CDNS_765158635885 $T=10820 5970 0 0 $X=10740 $Y=5840
X11 8 M2_M1_CDNS_765158635885 $T=11040 2940 0 0 $X=10960 $Y=2810
X12 2 M2_M1_CDNS_765158635885 $T=11390 3320 0 0 $X=11310 $Y=3190
X13 7 M2_M1_CDNS_765158635885 $T=12920 3510 0 0 $X=12840 $Y=3380
X14 4 M2_M1_CDNS_7651586358826 $T=6470 5920 0 0 $X=6340 $Y=5790
X15 3 M2_M1_CDNS_7651586358826 $T=7620 3360 0 0 $X=7490 $Y=3230
X16 3 M2_M1_CDNS_7651586358826 $T=10320 3640 0 0 $X=10190 $Y=3510
X17 4 M2_M1_CDNS_7651586358827 $T=3420 5920 0 0 $X=3290 $Y=5790
X18 10 4 7 5 inv $T=12350 3410 0 0 $X=11870 $Y=1250
X19 1 4 5 11 9 2 xor $T=4170 3810 0 0 $X=1950 $Y=1250
X20 9 4 5 8 6 3 xor $T=8070 3810 0 0 $X=5850 $Y=1250
X21 3 M3_M2_CDNS_7651586358835 $T=7300 3360 0 0 $X=7170 $Y=3230
X22 3 M3_M2_CDNS_7651586358835 $T=10110 3640 0 0 $X=9980 $Y=3510
X23 10 9 3 4 8 5 2 12 13 14
+ 15 fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 11 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 4 1 11 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 2 1 9 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 8 9 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 4 9 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 3 9 6 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 7 10 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 4 10 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pipeline_mult                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pipeline_mult 4 3 14 13 42 43 44 45 46 58
+ 57 56 59 60 61 62 63 47 2 1
** N=199 EP=20 FDC=697
X0 1 M10_M9_CDNS_765158635880 $T=17800 31890 0 0 $X=16840 $Y=31610
X1 1 M10_M9_CDNS_765158635880 $T=17800 41250 0 0 $X=16840 $Y=40970
X2 1 M10_M9_CDNS_765158635880 $T=17800 52810 0 0 $X=16840 $Y=52530
X3 1 M10_M9_CDNS_765158635880 $T=17800 62670 0 0 $X=16840 $Y=62390
X4 2 M10_M9_CDNS_765158635880 $T=19460 36430 0 0 $X=18500 $Y=36150
X5 2 M10_M9_CDNS_765158635880 $T=19460 42880 0 0 $X=18500 $Y=42600
X6 2 M10_M9_CDNS_765158635880 $T=19460 57580 0 0 $X=18500 $Y=57300
X7 2 M10_M9_CDNS_765158635880 $T=19970 67840 0 0 $X=19010 $Y=67560
X8 1 M10_M9_CDNS_765158635880 $T=25170 26020 0 0 $X=24210 $Y=25740
X9 1 M10_M9_CDNS_765158635880 $T=25170 36360 0 0 $X=24210 $Y=36080
X10 1 M10_M9_CDNS_765158635880 $T=26180 46200 0 0 $X=25220 $Y=45920
X11 1 M10_M9_CDNS_765158635880 $T=26180 55950 0 0 $X=25220 $Y=55670
X12 2 M10_M9_CDNS_765158635880 $T=29850 33170 0 0 $X=28890 $Y=32890
X13 2 M10_M9_CDNS_765158635880 $T=29850 41710 0 0 $X=28890 $Y=41430
X14 2 M10_M9_CDNS_765158635880 $T=29850 49920 0 0 $X=28890 $Y=49640
X15 2 M10_M9_CDNS_765158635880 $T=29850 60150 0 0 $X=28890 $Y=59870
X16 1 M10_M9_CDNS_765158635880 $T=31640 27280 0 0 $X=30680 $Y=27000
X17 1 M10_M9_CDNS_765158635880 $T=31640 36120 0 0 $X=30680 $Y=35840
X18 1 M10_M9_CDNS_765158635880 $T=31640 43460 0 0 $X=30680 $Y=43180
X19 1 M10_M9_CDNS_765158635880 $T=31640 51990 0 0 $X=30680 $Y=51710
X20 1 M10_M9_CDNS_765158635880 $T=47370 27000 0 0 $X=46410 $Y=26720
X21 1 M10_M9_CDNS_765158635880 $T=47370 34350 0 0 $X=46410 $Y=34070
X22 1 M10_M9_CDNS_765158635880 $T=48190 19140 0 0 $X=47230 $Y=18860
X23 1 M10_M9_CDNS_765158635880 $T=50320 1650 0 0 $X=49360 $Y=1370
X24 1 M10_M9_CDNS_765158635880 $T=50560 43090 0 0 $X=49600 $Y=42810
X25 2 M10_M9_CDNS_765158635880 $T=52000 24420 0 0 $X=51040 $Y=24140
X26 2 M10_M9_CDNS_765158635880 $T=52000 32940 0 0 $X=51040 $Y=32660
X27 2 M10_M9_CDNS_765158635880 $T=52000 41710 0 0 $X=51040 $Y=41430
X28 2 M10_M9_CDNS_765158635880 $T=52000 50750 0 0 $X=51040 $Y=50470
X29 2 M10_M9_CDNS_765158635880 $T=52000 70000 0 0 $X=51040 $Y=69720
X30 1 M10_M9_CDNS_765158635880 $T=54310 36140 0 0 $X=53350 $Y=35860
X31 1 M10_M9_CDNS_765158635880 $T=57590 19010 0 0 $X=56630 $Y=18730
X32 1 M10_M9_CDNS_765158635880 $T=57590 27220 0 0 $X=56630 $Y=26940
X33 1 M10_M9_CDNS_765158635880 $T=58810 43360 0 0 $X=57850 $Y=43080
X34 1 M10_M9_CDNS_765158635880 $T=74710 18390 0 0 $X=73750 $Y=18110
X35 1 M10_M9_CDNS_765158635880 $T=74710 26320 0 0 $X=73750 $Y=26040
X36 1 M10_M9_CDNS_765158635880 $T=74710 34190 0 0 $X=73750 $Y=33910
X37 1 M10_M9_CDNS_765158635880 $T=74880 9960 0 0 $X=73920 $Y=9680
X38 2 M10_M9_CDNS_765158635880 $T=77130 16720 0 0 $X=76170 $Y=16440
X39 2 M10_M9_CDNS_765158635880 $T=77130 24150 0 0 $X=76170 $Y=23870
X40 2 M10_M9_CDNS_765158635880 $T=77130 33380 0 0 $X=76170 $Y=33100
X41 2 M10_M9_CDNS_765158635880 $T=78960 40520 0 0 $X=78000 $Y=40240
X42 1 M10_M9_CDNS_765158635880 $T=83500 11210 0 0 $X=82540 $Y=10930
X43 1 M10_M9_CDNS_765158635880 $T=85120 19060 0 0 $X=84160 $Y=18780
X44 1 M10_M9_CDNS_765158635880 $T=85120 28410 0 0 $X=84160 $Y=28130
X45 1 M10_M9_CDNS_765158635880 $T=85120 35190 0 0 $X=84160 $Y=34910
X46 2 M10_M9_CDNS_765158635880 $T=99950 62120 0 0 $X=98990 $Y=61840
X47 2 M10_M9_CDNS_765158635880 $T=100620 51980 0 0 $X=99660 $Y=51700
X48 2 M10_M9_CDNS_765158635880 $T=102130 14020 0 0 $X=101170 $Y=13740
X49 2 M10_M9_CDNS_765158635880 $T=102130 22060 0 0 $X=101170 $Y=21780
X50 2 M10_M9_CDNS_765158635880 $T=102130 29250 0 0 $X=101170 $Y=28970
X51 2 M10_M9_CDNS_765158635880 $T=102130 38320 0 0 $X=101170 $Y=38040
X52 2 M10_M9_CDNS_765158635880 $T=105780 67340 0 0 $X=104820 $Y=67060
X53 1 M10_M9_CDNS_765158635880 $T=106700 9960 0 0 $X=105740 $Y=9680
X54 1 M10_M9_CDNS_765158635880 $T=106700 18350 0 0 $X=105740 $Y=18070
X55 1 M10_M9_CDNS_765158635880 $T=106700 26740 0 0 $X=105740 $Y=26460
X56 1 M10_M9_CDNS_765158635880 $T=106700 35130 0 0 $X=105740 $Y=34850
X57 1 M10_M9_CDNS_765158635880 $T=106700 46110 0 0 $X=105740 $Y=45830
X58 1 M10_M9_CDNS_765158635880 $T=106700 55990 0 0 $X=105740 $Y=55710
X59 1 M10_M9_CDNS_765158635880 $T=106700 61440 0 0 $X=105740 $Y=61160
X60 3 M4_M3_CDNS_765158635881 $T=10310 56470 0 0 $X=9870 $Y=56060
X61 4 M4_M3_CDNS_765158635881 $T=10500 65720 0 0 $X=10060 $Y=65310
X62 5 M4_M3_CDNS_765158635882 $T=44180 28360 0 0 $X=44100 $Y=28230
X63 6 M4_M3_CDNS_765158635882 $T=44940 37650 0 0 $X=44860 $Y=37520
X64 7 M4_M3_CDNS_765158635882 $T=46460 45180 0 0 $X=46380 $Y=45050
X65 8 M4_M3_CDNS_765158635882 $T=47910 54210 0 0 $X=47830 $Y=54080
X66 5 M4_M3_CDNS_765158635882 $T=48980 28360 0 0 $X=48900 $Y=28230
X67 6 M4_M3_CDNS_765158635882 $T=49760 37640 0 0 $X=49680 $Y=37510
X68 7 M4_M3_CDNS_765158635882 $T=52850 45180 0 0 $X=52770 $Y=45050
X69 9 M4_M3_CDNS_765158635882 $T=70440 19260 0 0 $X=70360 $Y=19130
X70 10 M4_M3_CDNS_765158635882 $T=70650 27640 0 0 $X=70570 $Y=27510
X71 11 M4_M3_CDNS_765158635882 $T=71540 35870 0 0 $X=71460 $Y=35740
X72 12 M4_M3_CDNS_765158635882 $T=72680 45660 0 0 $X=72600 $Y=45530
X73 9 M4_M3_CDNS_765158635882 $T=74880 19260 0 0 $X=74800 $Y=19130
X74 10 M4_M3_CDNS_765158635882 $T=76020 27640 0 0 $X=75940 $Y=27510
X75 11 M4_M3_CDNS_765158635882 $T=76960 35860 0 0 $X=76880 $Y=35730
X76 12 M4_M3_CDNS_765158635882 $T=96080 50090 0 0 $X=96000 $Y=49960
X77 8 M4_M3_CDNS_765158635882 $T=96940 60090 0 0 $X=96860 $Y=59960
X78 13 M4_M3_CDNS_765158635883 $T=10290 35240 0 0 $X=9930 $Y=34750
X79 14 M4_M3_CDNS_765158635883 $T=10390 44020 0 0 $X=10030 $Y=43530
X80 15 M3_M2_CDNS_765158635884 $T=25130 29430 0 0 $X=25050 $Y=29300
X81 16 M3_M2_CDNS_765158635884 $T=28320 39590 0 0 $X=28240 $Y=39460
X82 17 M3_M2_CDNS_765158635884 $T=28520 47670 0 0 $X=28440 $Y=47540
X83 18 M3_M2_CDNS_765158635884 $T=28930 38580 0 0 $X=28850 $Y=38450
X84 19 M3_M2_CDNS_765158635884 $T=28970 37640 0 0 $X=28890 $Y=37510
X85 20 M3_M2_CDNS_765158635884 $T=29860 45980 0 0 $X=29780 $Y=45850
X86 21 M3_M2_CDNS_765158635884 $T=29870 46920 0 0 $X=29790 $Y=46790
X87 22 M3_M2_CDNS_765158635884 $T=31070 31220 0 0 $X=30990 $Y=31090
X88 23 M3_M2_CDNS_765158635884 $T=32300 55080 0 0 $X=32220 $Y=54950
X89 24 M3_M2_CDNS_765158635884 $T=32310 54610 0 0 $X=32230 $Y=54480
X90 25 M3_M2_CDNS_765158635884 $T=49150 30450 0 0 $X=49070 $Y=30320
X91 26 M3_M2_CDNS_765158635884 $T=49160 21810 0 0 $X=49080 $Y=21680
X92 27 M3_M2_CDNS_765158635884 $T=50340 21230 0 0 $X=50260 $Y=21100
X93 28 M3_M2_CDNS_765158635884 $T=51060 38580 0 0 $X=50980 $Y=38450
X94 29 M3_M2_CDNS_765158635884 $T=52900 46770 0 0 $X=52820 $Y=46640
X95 30 M3_M2_CDNS_765158635884 $T=53940 29990 0 0 $X=53860 $Y=29860
X96 31 M3_M2_CDNS_765158635884 $T=54020 38140 0 0 $X=53940 $Y=38010
X97 32 M3_M2_CDNS_765158635884 $T=54070 21740 0 0 $X=53990 $Y=21610
X98 33 M3_M2_CDNS_765158635884 $T=75930 21540 0 0 $X=75850 $Y=21410
X99 34 M3_M2_CDNS_765158635884 $T=76120 13000 0 0 $X=76040 $Y=12870
X100 35 M3_M2_CDNS_765158635884 $T=76270 29940 0 0 $X=76190 $Y=29810
X101 34 M3_M2_CDNS_765158635884 $T=83280 16240 0 0 $X=83200 $Y=16110
X102 33 M3_M2_CDNS_765158635884 $T=83280 23710 0 0 $X=83200 $Y=23580
X103 35 M3_M2_CDNS_765158635884 $T=83280 32890 0 0 $X=83200 $Y=32760
X104 9 M3_M2_CDNS_765158635884 $T=92880 19820 0 0 $X=92800 $Y=19690
X105 10 M3_M2_CDNS_765158635884 $T=92880 29000 0 0 $X=92800 $Y=28870
X106 11 M3_M2_CDNS_765158635884 $T=92880 36230 0 0 $X=92800 $Y=36100
X107 12 M3_M2_CDNS_765158635884 $T=99140 50130 0 0 $X=99060 $Y=50000
X108 8 M3_M2_CDNS_765158635884 $T=99140 60130 0 0 $X=99060 $Y=60000
X109 36 M3_M2_CDNS_765158635884 $T=104800 29590 0 0 $X=104720 $Y=29460
X110 37 M3_M2_CDNS_765158635884 $T=104890 12740 0 0 $X=104810 $Y=12610
X111 38 M3_M2_CDNS_765158635884 $T=105170 21180 0 0 $X=105090 $Y=21050
X112 24 M2_M1_CDNS_765158635885 $T=16610 55790 0 0 $X=16530 $Y=55660
X113 39 M2_M1_CDNS_765158635885 $T=16620 65580 0 0 $X=16540 $Y=65450
X114 19 M2_M1_CDNS_765158635885 $T=16910 35060 0 0 $X=16830 $Y=34930
X115 20 M2_M1_CDNS_765158635885 $T=16910 44530 0 0 $X=16830 $Y=44400
X116 15 M2_M1_CDNS_765158635885 $T=25130 29430 0 0 $X=25050 $Y=29300
X117 21 M2_M1_CDNS_765158635885 $T=25230 48920 0 0 $X=25150 $Y=48790
X118 23 M2_M1_CDNS_765158635885 $T=25230 58750 0 0 $X=25150 $Y=58620
X119 18 M2_M1_CDNS_765158635885 $T=25240 39680 0 0 $X=25160 $Y=39550
X120 26 M2_M1_CDNS_765158635885 $T=46750 21820 0 0 $X=46670 $Y=21690
X121 25 M2_M1_CDNS_765158635885 $T=47610 30450 0 0 $X=47530 $Y=30320
X122 28 M2_M1_CDNS_765158635885 $T=48850 38580 0 0 $X=48770 $Y=38450
X123 29 M2_M1_CDNS_765158635885 $T=50700 46770 0 0 $X=50620 $Y=46640
X124 34 M2_M1_CDNS_765158635885 $T=73180 12220 0 0 $X=73100 $Y=12090
X125 33 M2_M1_CDNS_765158635885 $T=73440 21500 0 0 $X=73360 $Y=21370
X126 35 M2_M1_CDNS_765158635885 $T=73980 29570 0 0 $X=73900 $Y=29440
X127 40 M2_M1_CDNS_765158635885 $T=75410 37650 0 0 $X=75330 $Y=37520
X128 34 M2_M1_CDNS_765158635885 $T=84630 16240 0 0 $X=84550 $Y=16110
X129 33 M2_M1_CDNS_765158635885 $T=84630 23710 0 0 $X=84550 $Y=23580
X130 35 M2_M1_CDNS_765158635885 $T=84630 32890 0 0 $X=84550 $Y=32760
X131 40 M2_M1_CDNS_765158635885 $T=84630 40120 0 0 $X=84550 $Y=39990
X132 41 M2_M1_CDNS_765158635885 $T=94230 12350 0 0 $X=94150 $Y=12220
X133 9 M2_M1_CDNS_765158635885 $T=94230 19820 0 0 $X=94150 $Y=19690
X134 10 M2_M1_CDNS_765158635885 $T=94230 29000 0 0 $X=94150 $Y=28870
X135 11 M2_M1_CDNS_765158635885 $T=94230 36230 0 0 $X=94150 $Y=36100
X136 12 M2_M1_CDNS_765158635885 $T=100490 50130 0 0 $X=100410 $Y=50000
X137 8 M2_M1_CDNS_765158635885 $T=100490 60130 0 0 $X=100410 $Y=60000
X138 39 M2_M1_CDNS_765158635885 $T=105900 65540 0 0 $X=105820 $Y=65410
X139 3 M4_M3_CDNS_765158635886 $T=13300 55730 0 0 $X=13220 $Y=55320
X140 4 M4_M3_CDNS_765158635886 $T=13300 65530 0 0 $X=13220 $Y=65120
X141 13 M4_M3_CDNS_765158635886 $T=13600 35000 0 0 $X=13520 $Y=34590
X142 14 M4_M3_CDNS_765158635886 $T=13600 44460 0 0 $X=13520 $Y=44050
X143 13 M4_M3_CDNS_765158635886 $T=21820 29380 0 0 $X=21740 $Y=28970
X144 4 M4_M3_CDNS_765158635886 $T=21910 58670 0 0 $X=21830 $Y=58260
X145 14 M4_M3_CDNS_765158635886 $T=21920 39620 0 0 $X=21840 $Y=39210
X146 3 M4_M3_CDNS_765158635886 $T=21920 48870 0 0 $X=21840 $Y=48460
X147 13 M4_M3_CDNS_765158635886 $T=43440 21760 0 0 $X=43360 $Y=21350
X148 14 M4_M3_CDNS_765158635886 $T=44290 30400 0 0 $X=44210 $Y=29990
X149 3 M4_M3_CDNS_765158635886 $T=45490 38520 0 0 $X=45410 $Y=38110
X150 4 M4_M3_CDNS_765158635886 $T=47380 46710 0 0 $X=47300 $Y=46300
X151 13 M4_M3_CDNS_765158635886 $T=69880 12180 0 0 $X=69800 $Y=11770
X152 14 M4_M3_CDNS_765158635886 $T=70120 21430 0 0 $X=70040 $Y=21020
X153 3 M4_M3_CDNS_765158635886 $T=70670 29530 0 0 $X=70590 $Y=29120
X154 4 M4_M3_CDNS_765158635886 $T=72100 37590 0 0 $X=72020 $Y=37180
X155 3 M2_M1_CDNS_765158635887 $T=13300 55730 0 0 $X=13220 $Y=55320
X156 4 M2_M1_CDNS_765158635887 $T=13300 65530 0 0 $X=13220 $Y=65120
X157 13 M2_M1_CDNS_765158635887 $T=13600 35000 0 0 $X=13520 $Y=34590
X158 14 M2_M1_CDNS_765158635887 $T=13600 44460 0 0 $X=13520 $Y=44050
X159 42 M2_M1_CDNS_765158635887 $T=14600 55440 0 0 $X=14520 $Y=55030
X160 42 M2_M1_CDNS_765158635887 $T=14600 65230 0 0 $X=14520 $Y=64820
X161 42 M2_M1_CDNS_765158635887 $T=14900 34700 0 0 $X=14820 $Y=34290
X162 42 M2_M1_CDNS_765158635887 $T=14900 44170 0 0 $X=14820 $Y=43760
X163 13 M2_M1_CDNS_765158635887 $T=21820 29380 0 0 $X=21740 $Y=28970
X164 14 M2_M1_CDNS_765158635887 $T=21920 39620 0 0 $X=21840 $Y=39210
X165 3 M2_M1_CDNS_765158635887 $T=21920 48870 0 0 $X=21840 $Y=48460
X166 4 M2_M1_CDNS_765158635887 $T=21920 58680 0 0 $X=21840 $Y=58270
X167 43 M2_M1_CDNS_765158635887 $T=23120 29070 0 0 $X=23040 $Y=28660
X168 43 M2_M1_CDNS_765158635887 $T=23220 39320 0 0 $X=23140 $Y=38910
X169 43 M2_M1_CDNS_765158635887 $T=23220 48570 0 0 $X=23140 $Y=48160
X170 43 M2_M1_CDNS_765158635887 $T=23220 58400 0 0 $X=23140 $Y=57990
X171 13 M2_M1_CDNS_765158635887 $T=43440 21760 0 0 $X=43360 $Y=21350
X172 14 M2_M1_CDNS_765158635887 $T=44290 30400 0 0 $X=44210 $Y=29990
X173 44 M2_M1_CDNS_765158635887 $T=44740 21460 0 0 $X=44660 $Y=21050
X174 3 M2_M1_CDNS_765158635887 $T=45490 38520 0 0 $X=45410 $Y=38110
X175 44 M2_M1_CDNS_765158635887 $T=45590 30100 0 0 $X=45510 $Y=29690
X176 44 M2_M1_CDNS_765158635887 $T=46790 38220 0 0 $X=46710 $Y=37810
X177 4 M2_M1_CDNS_765158635887 $T=47380 46710 0 0 $X=47300 $Y=46300
X178 44 M2_M1_CDNS_765158635887 $T=48680 46410 0 0 $X=48600 $Y=46000
X179 13 M2_M1_CDNS_765158635887 $T=69880 12180 0 0 $X=69800 $Y=11770
X180 14 M2_M1_CDNS_765158635887 $T=70120 21430 0 0 $X=70040 $Y=21020
X181 3 M2_M1_CDNS_765158635887 $T=70670 29530 0 0 $X=70590 $Y=29120
X182 45 M2_M1_CDNS_765158635887 $T=71180 11870 0 0 $X=71100 $Y=11460
X183 45 M2_M1_CDNS_765158635887 $T=71420 21130 0 0 $X=71340 $Y=20720
X184 45 M2_M1_CDNS_765158635887 $T=71970 29230 0 0 $X=71890 $Y=28820
X185 4 M2_M1_CDNS_765158635887 $T=72100 37590 0 0 $X=72020 $Y=37180
X186 45 M2_M1_CDNS_765158635887 $T=73400 37290 0 0 $X=73320 $Y=36880
X187 3 M3_M2_CDNS_765158635888 $T=13300 55730 0 0 $X=13220 $Y=55320
X188 4 M3_M2_CDNS_765158635888 $T=13300 65530 0 0 $X=13220 $Y=65120
X189 13 M3_M2_CDNS_765158635888 $T=13600 35000 0 0 $X=13520 $Y=34590
X190 14 M3_M2_CDNS_765158635888 $T=13600 44460 0 0 $X=13520 $Y=44050
X191 42 M3_M2_CDNS_765158635888 $T=14600 55440 0 0 $X=14520 $Y=55030
X192 42 M3_M2_CDNS_765158635888 $T=14600 65230 0 0 $X=14520 $Y=64820
X193 42 M3_M2_CDNS_765158635888 $T=14900 34700 0 0 $X=14820 $Y=34290
X194 42 M3_M2_CDNS_765158635888 $T=14900 44170 0 0 $X=14820 $Y=43760
X195 13 M3_M2_CDNS_765158635888 $T=21820 29380 0 0 $X=21740 $Y=28970
X196 14 M3_M2_CDNS_765158635888 $T=21920 39620 0 0 $X=21840 $Y=39210
X197 3 M3_M2_CDNS_765158635888 $T=21920 48870 0 0 $X=21840 $Y=48460
X198 4 M3_M2_CDNS_765158635888 $T=21920 58680 0 0 $X=21840 $Y=58270
X199 43 M3_M2_CDNS_765158635888 $T=23120 29070 0 0 $X=23040 $Y=28660
X200 43 M3_M2_CDNS_765158635888 $T=23220 39320 0 0 $X=23140 $Y=38910
X201 43 M3_M2_CDNS_765158635888 $T=23220 48570 0 0 $X=23140 $Y=48160
X202 43 M3_M2_CDNS_765158635888 $T=23220 58400 0 0 $X=23140 $Y=57990
X203 13 M3_M2_CDNS_765158635888 $T=43440 21760 0 0 $X=43360 $Y=21350
X204 14 M3_M2_CDNS_765158635888 $T=44290 30400 0 0 $X=44210 $Y=29990
X205 44 M3_M2_CDNS_765158635888 $T=44740 21460 0 0 $X=44660 $Y=21050
X206 3 M3_M2_CDNS_765158635888 $T=45490 38520 0 0 $X=45410 $Y=38110
X207 44 M3_M2_CDNS_765158635888 $T=45590 30100 0 0 $X=45510 $Y=29690
X208 44 M3_M2_CDNS_765158635888 $T=46790 38220 0 0 $X=46710 $Y=37810
X209 4 M3_M2_CDNS_765158635888 $T=47380 46710 0 0 $X=47300 $Y=46300
X210 44 M3_M2_CDNS_765158635888 $T=48680 46410 0 0 $X=48600 $Y=46000
X211 13 M3_M2_CDNS_765158635888 $T=69880 12180 0 0 $X=69800 $Y=11770
X212 14 M3_M2_CDNS_765158635888 $T=70120 21430 0 0 $X=70040 $Y=21020
X213 3 M3_M2_CDNS_765158635888 $T=70670 29530 0 0 $X=70590 $Y=29120
X214 45 M3_M2_CDNS_765158635888 $T=71180 11870 0 0 $X=71100 $Y=11460
X215 45 M3_M2_CDNS_765158635888 $T=71420 21130 0 0 $X=71340 $Y=20720
X216 45 M3_M2_CDNS_765158635888 $T=71970 29230 0 0 $X=71890 $Y=28820
X217 4 M3_M2_CDNS_765158635888 $T=72100 37590 0 0 $X=72020 $Y=37180
X218 45 M3_M2_CDNS_765158635888 $T=73400 37290 0 0 $X=73320 $Y=36880
X219 46 M4_M3_CDNS_765158635889 $T=83660 22300 0 0 $X=83440 $Y=22170
X220 46 M4_M3_CDNS_765158635889 $T=83660 31480 0 0 $X=83440 $Y=31350
X221 46 M4_M3_CDNS_765158635889 $T=83660 38710 0 0 $X=83440 $Y=38580
X222 46 M4_M3_CDNS_765158635889 $T=83670 14830 0 0 $X=83450 $Y=14700
X223 47 M4_M3_CDNS_765158635889 $T=91230 14480 0 0 $X=91010 $Y=14350
X224 47 M4_M3_CDNS_765158635889 $T=91230 21950 0 0 $X=91010 $Y=21820
X225 47 M4_M3_CDNS_765158635889 $T=91230 31130 0 0 $X=91010 $Y=31000
X226 47 M4_M3_CDNS_765158635889 $T=91230 38320 0 0 $X=91010 $Y=38190
X227 46 M4_M3_CDNS_765158635889 $T=93250 42620 0 0 $X=93030 $Y=42490
X228 46 M4_M3_CDNS_765158635889 $T=93250 44610 0 0 $X=93030 $Y=44480
X229 46 M4_M3_CDNS_765158635889 $T=93260 10940 0 0 $X=93040 $Y=10810
X230 46 M4_M3_CDNS_765158635889 $T=93260 18410 0 0 $X=93040 $Y=18280
X231 46 M4_M3_CDNS_765158635889 $T=93260 27590 0 0 $X=93040 $Y=27460
X232 46 M4_M3_CDNS_765158635889 $T=93260 34820 0 0 $X=93040 $Y=34690
X233 46 M4_M3_CDNS_765158635889 $T=99510 58720 0 0 $X=99290 $Y=58590
X234 46 M4_M3_CDNS_765158635889 $T=99520 48720 0 0 $X=99300 $Y=48590
X235 47 M4_M3_CDNS_765158635889 $T=100830 10590 0 180 $X=100610 $Y=10460
X236 47 M4_M3_CDNS_765158635889 $T=100830 18060 0 180 $X=100610 $Y=17930
X237 47 M4_M3_CDNS_765158635889 $T=100830 27240 0 180 $X=100610 $Y=27110
X238 47 M4_M3_CDNS_765158635889 $T=100830 34470 0 0 $X=100610 $Y=34340
X239 46 M4_M3_CDNS_765158635889 $T=101070 68620 0 0 $X=100850 $Y=68490
X240 46 M4_M3_CDNS_765158635889 $T=104930 64130 0 0 $X=104710 $Y=64000
X241 47 M4_M3_CDNS_765158635889 $T=107050 58360 0 0 $X=106830 $Y=58230
X242 47 M4_M3_CDNS_765158635889 $T=107080 48320 0 0 $X=106860 $Y=48190
X243 47 M4_M3_CDNS_765158635889 $T=112490 63750 0 0 $X=112270 $Y=63620
X244 47 M4_M3_CDNS_765158635889 $T=112490 68450 0 0 $X=112270 $Y=68320
X245 2 M11_M10_CDNS_7651586358810 $T=19460 36430 0 0 $X=18500 $Y=36150
X246 2 M11_M10_CDNS_7651586358810 $T=19460 42880 0 0 $X=18500 $Y=42600
X247 2 M11_M10_CDNS_7651586358810 $T=19460 57580 0 0 $X=18500 $Y=57300
X248 2 M11_M10_CDNS_7651586358810 $T=19970 67840 0 0 $X=19010 $Y=67560
X249 2 M11_M10_CDNS_7651586358810 $T=29850 33170 0 0 $X=28890 $Y=32890
X250 2 M11_M10_CDNS_7651586358810 $T=29850 41710 0 0 $X=28890 $Y=41430
X251 2 M11_M10_CDNS_7651586358810 $T=29850 49920 0 0 $X=28890 $Y=49640
X252 2 M11_M10_CDNS_7651586358810 $T=29850 60150 0 0 $X=28890 $Y=59870
X253 1 M11_M10_CDNS_7651586358810 $T=50320 1650 0 0 $X=49360 $Y=1370
X254 2 M11_M10_CDNS_7651586358810 $T=52000 24420 0 0 $X=51040 $Y=24140
X255 2 M11_M10_CDNS_7651586358810 $T=52000 32940 0 0 $X=51040 $Y=32660
X256 2 M11_M10_CDNS_7651586358810 $T=52000 41710 0 0 $X=51040 $Y=41430
X257 2 M11_M10_CDNS_7651586358810 $T=52000 50750 0 0 $X=51040 $Y=50470
X258 2 M11_M10_CDNS_7651586358810 $T=52000 70000 0 0 $X=51040 $Y=69720
X259 2 M11_M10_CDNS_7651586358810 $T=77130 16720 0 0 $X=76170 $Y=16440
X260 2 M11_M10_CDNS_7651586358810 $T=77130 24150 0 0 $X=76170 $Y=23870
X261 2 M11_M10_CDNS_7651586358810 $T=77130 33380 0 0 $X=76170 $Y=33100
X262 2 M11_M10_CDNS_7651586358810 $T=78960 40520 0 0 $X=78000 $Y=40240
X263 2 M11_M10_CDNS_7651586358810 $T=99950 62120 0 0 $X=98990 $Y=61840
X264 2 M11_M10_CDNS_7651586358810 $T=100620 51980 0 0 $X=99660 $Y=51700
X265 2 M11_M10_CDNS_7651586358810 $T=102130 14020 0 0 $X=101170 $Y=13740
X266 2 M11_M10_CDNS_7651586358810 $T=102130 22060 0 0 $X=101170 $Y=21780
X267 2 M11_M10_CDNS_7651586358810 $T=102130 29250 0 0 $X=101170 $Y=28970
X268 2 M11_M10_CDNS_7651586358810 $T=102130 38320 0 0 $X=101170 $Y=38040
X269 2 M11_M10_CDNS_7651586358810 $T=105780 67340 0 0 $X=104820 $Y=67060
X270 13 M5_M4_CDNS_7651586358811 $T=43590 35230 0 0 $X=43510 $Y=35100
X271 14 M5_M4_CDNS_7651586358811 $T=44450 44030 0 0 $X=44370 $Y=43900
X272 13 M5_M4_CDNS_7651586358811 $T=44970 35230 0 0 $X=44890 $Y=35100
X273 3 M5_M4_CDNS_7651586358811 $T=45820 56470 0 0 $X=45740 $Y=56340
X274 14 M5_M4_CDNS_7651586358811 $T=46380 44030 0 0 $X=46300 $Y=43900
X275 3 M5_M4_CDNS_7651586358811 $T=49010 56470 0 0 $X=48930 $Y=56340
X276 8 M5_M4_CDNS_7651586358811 $T=69610 54210 0 0 $X=69530 $Y=54080
X277 8 M5_M4_CDNS_7651586358811 $T=74290 54220 0 0 $X=74210 $Y=54090
X278 1 M5_M4_CDNS_7651586358812 $T=17800 31900 0 0 $X=17440 $Y=31770
X279 1 M5_M4_CDNS_7651586358812 $T=17800 41260 0 0 $X=17440 $Y=41130
X280 1 M5_M4_CDNS_7651586358812 $T=17800 52820 0 0 $X=17440 $Y=52690
X281 1 M5_M4_CDNS_7651586358812 $T=17800 62680 0 0 $X=17440 $Y=62550
X282 2 M5_M4_CDNS_7651586358812 $T=19460 36430 0 0 $X=19100 $Y=36300
X283 2 M5_M4_CDNS_7651586358812 $T=19460 42880 0 0 $X=19100 $Y=42750
X284 2 M5_M4_CDNS_7651586358812 $T=19460 57580 0 0 $X=19100 $Y=57450
X285 2 M5_M4_CDNS_7651586358812 $T=19970 67840 0 0 $X=19610 $Y=67710
X286 1 M5_M4_CDNS_7651586358812 $T=25170 26030 0 0 $X=24810 $Y=25900
X287 1 M5_M4_CDNS_7651586358812 $T=25170 36370 0 0 $X=24810 $Y=36240
X288 1 M5_M4_CDNS_7651586358812 $T=26180 46210 0 0 $X=25820 $Y=46080
X289 1 M5_M4_CDNS_7651586358812 $T=26180 55960 0 0 $X=25820 $Y=55830
X290 2 M5_M4_CDNS_7651586358812 $T=29850 33170 0 0 $X=29490 $Y=33040
X291 2 M5_M4_CDNS_7651586358812 $T=29850 41710 0 0 $X=29490 $Y=41580
X292 2 M5_M4_CDNS_7651586358812 $T=29850 49920 0 0 $X=29490 $Y=49790
X293 2 M5_M4_CDNS_7651586358812 $T=29850 60150 0 0 $X=29490 $Y=60020
X294 1 M5_M4_CDNS_7651586358812 $T=31640 27290 0 0 $X=31280 $Y=27160
X295 1 M5_M4_CDNS_7651586358812 $T=31640 36130 0 0 $X=31280 $Y=36000
X296 1 M5_M4_CDNS_7651586358812 $T=31640 43470 0 0 $X=31280 $Y=43340
X297 1 M5_M4_CDNS_7651586358812 $T=31640 52000 0 0 $X=31280 $Y=51870
X298 1 M5_M4_CDNS_7651586358812 $T=47370 27010 0 0 $X=47010 $Y=26880
X299 1 M5_M4_CDNS_7651586358812 $T=47370 34360 0 0 $X=47010 $Y=34230
X300 1 M5_M4_CDNS_7651586358812 $T=48190 19140 0 0 $X=47830 $Y=19010
X301 1 M5_M4_CDNS_7651586358812 $T=50630 43060 0 0 $X=50270 $Y=42930
X302 2 M5_M4_CDNS_7651586358812 $T=52000 24420 0 0 $X=51640 $Y=24290
X303 2 M5_M4_CDNS_7651586358812 $T=52000 32940 0 0 $X=51640 $Y=32810
X304 2 M5_M4_CDNS_7651586358812 $T=52000 41710 0 0 $X=51640 $Y=41580
X305 2 M5_M4_CDNS_7651586358812 $T=52000 50750 0 0 $X=51640 $Y=50620
X306 2 M5_M4_CDNS_7651586358812 $T=52000 70000 0 0 $X=51640 $Y=69870
X307 1 M5_M4_CDNS_7651586358812 $T=54300 36130 0 0 $X=53940 $Y=36000
X308 1 M5_M4_CDNS_7651586358812 $T=57590 18970 0 0 $X=57230 $Y=18840
X309 1 M5_M4_CDNS_7651586358812 $T=57590 27180 0 0 $X=57230 $Y=27050
X310 1 M5_M4_CDNS_7651586358812 $T=58810 43370 0 0 $X=58450 $Y=43240
X311 1 M5_M4_CDNS_7651586358812 $T=74710 18350 0 0 $X=74350 $Y=18220
X312 1 M5_M4_CDNS_7651586358812 $T=74710 26280 0 0 $X=74350 $Y=26150
X313 1 M5_M4_CDNS_7651586358812 $T=74710 34150 0 0 $X=74350 $Y=34020
X314 1 M5_M4_CDNS_7651586358812 $T=74880 9920 0 0 $X=74520 $Y=9790
X315 2 M5_M4_CDNS_7651586358812 $T=77130 16720 0 0 $X=76770 $Y=16590
X316 2 M5_M4_CDNS_7651586358812 $T=77130 24150 0 0 $X=76770 $Y=24020
X317 2 M5_M4_CDNS_7651586358812 $T=77130 33380 0 0 $X=76770 $Y=33250
X318 2 M5_M4_CDNS_7651586358812 $T=78960 40520 0 0 $X=78600 $Y=40390
X319 1 M5_M4_CDNS_7651586358812 $T=83500 11170 0 0 $X=83140 $Y=11040
X320 1 M5_M4_CDNS_7651586358812 $T=85120 19020 0 0 $X=84760 $Y=18890
X321 1 M5_M4_CDNS_7651586358812 $T=85120 28370 0 0 $X=84760 $Y=28240
X322 1 M5_M4_CDNS_7651586358812 $T=85120 35150 0 0 $X=84760 $Y=35020
X323 2 M5_M4_CDNS_7651586358812 $T=99950 62120 0 0 $X=99590 $Y=61990
X324 2 M5_M4_CDNS_7651586358812 $T=100620 51980 0 0 $X=100260 $Y=51850
X325 2 M5_M4_CDNS_7651586358812 $T=102130 14020 0 0 $X=101770 $Y=13890
X326 2 M5_M4_CDNS_7651586358812 $T=102130 22060 0 0 $X=101770 $Y=21930
X327 2 M5_M4_CDNS_7651586358812 $T=102130 29250 0 0 $X=101770 $Y=29120
X328 2 M5_M4_CDNS_7651586358812 $T=102130 38320 0 0 $X=101770 $Y=38190
X329 2 M5_M4_CDNS_7651586358812 $T=105780 67340 0 0 $X=105420 $Y=67210
X330 1 M5_M4_CDNS_7651586358812 $T=106700 9920 0 0 $X=106340 $Y=9790
X331 1 M5_M4_CDNS_7651586358812 $T=106700 18310 0 0 $X=106340 $Y=18180
X332 1 M5_M4_CDNS_7651586358812 $T=106700 26700 0 0 $X=106340 $Y=26570
X333 1 M5_M4_CDNS_7651586358812 $T=106700 35090 0 0 $X=106340 $Y=34960
X334 1 M5_M4_CDNS_7651586358812 $T=106700 46070 0 0 $X=106340 $Y=45940
X335 1 M5_M4_CDNS_7651586358812 $T=106700 55950 0 0 $X=106340 $Y=55820
X336 1 M5_M4_CDNS_7651586358812 $T=106700 61400 0 0 $X=106340 $Y=61270
X337 1 M7_M6_CDNS_7651586358813 $T=17800 31900 0 0 $X=17440 $Y=31770
X338 1 M7_M6_CDNS_7651586358813 $T=17800 41260 0 0 $X=17440 $Y=41130
X339 1 M7_M6_CDNS_7651586358813 $T=17800 52820 0 0 $X=17440 $Y=52690
X340 1 M7_M6_CDNS_7651586358813 $T=17800 62680 0 0 $X=17440 $Y=62550
X341 2 M7_M6_CDNS_7651586358813 $T=19460 36430 0 0 $X=19100 $Y=36300
X342 2 M7_M6_CDNS_7651586358813 $T=19460 42880 0 0 $X=19100 $Y=42750
X343 2 M7_M6_CDNS_7651586358813 $T=19460 57580 0 0 $X=19100 $Y=57450
X344 2 M7_M6_CDNS_7651586358813 $T=19970 67840 0 0 $X=19610 $Y=67710
X345 1 M7_M6_CDNS_7651586358813 $T=25170 26030 0 0 $X=24810 $Y=25900
X346 1 M7_M6_CDNS_7651586358813 $T=25170 36370 0 0 $X=24810 $Y=36240
X347 1 M7_M6_CDNS_7651586358813 $T=26180 46210 0 0 $X=25820 $Y=46080
X348 1 M7_M6_CDNS_7651586358813 $T=26180 55960 0 0 $X=25820 $Y=55830
X349 2 M7_M6_CDNS_7651586358813 $T=29850 33170 0 0 $X=29490 $Y=33040
X350 2 M7_M6_CDNS_7651586358813 $T=29850 41710 0 0 $X=29490 $Y=41580
X351 2 M7_M6_CDNS_7651586358813 $T=29850 49920 0 0 $X=29490 $Y=49790
X352 2 M7_M6_CDNS_7651586358813 $T=29850 60150 0 0 $X=29490 $Y=60020
X353 1 M7_M6_CDNS_7651586358813 $T=31640 27290 0 0 $X=31280 $Y=27160
X354 1 M7_M6_CDNS_7651586358813 $T=31640 36130 0 0 $X=31280 $Y=36000
X355 1 M7_M6_CDNS_7651586358813 $T=31640 43470 0 0 $X=31280 $Y=43340
X356 1 M7_M6_CDNS_7651586358813 $T=31640 52000 0 0 $X=31280 $Y=51870
X357 1 M7_M6_CDNS_7651586358813 $T=47370 27010 0 0 $X=47010 $Y=26880
X358 1 M7_M6_CDNS_7651586358813 $T=47370 34360 0 0 $X=47010 $Y=34230
X359 1 M7_M6_CDNS_7651586358813 $T=48190 19140 0 0 $X=47830 $Y=19010
X360 1 M7_M6_CDNS_7651586358813 $T=50630 43060 0 0 $X=50270 $Y=42930
X361 2 M7_M6_CDNS_7651586358813 $T=52000 24420 0 0 $X=51640 $Y=24290
X362 2 M7_M6_CDNS_7651586358813 $T=52000 32940 0 0 $X=51640 $Y=32810
X363 2 M7_M6_CDNS_7651586358813 $T=52000 41710 0 0 $X=51640 $Y=41580
X364 2 M7_M6_CDNS_7651586358813 $T=52000 50750 0 0 $X=51640 $Y=50620
X365 2 M7_M6_CDNS_7651586358813 $T=52000 70000 0 0 $X=51640 $Y=69870
X366 1 M7_M6_CDNS_7651586358813 $T=54300 36130 0 0 $X=53940 $Y=36000
X367 1 M7_M6_CDNS_7651586358813 $T=57590 18970 0 0 $X=57230 $Y=18840
X368 1 M7_M6_CDNS_7651586358813 $T=57590 27180 0 0 $X=57230 $Y=27050
X369 1 M7_M6_CDNS_7651586358813 $T=58810 43370 0 0 $X=58450 $Y=43240
X370 1 M7_M6_CDNS_7651586358813 $T=74710 18350 0 0 $X=74350 $Y=18220
X371 1 M7_M6_CDNS_7651586358813 $T=74710 26280 0 0 $X=74350 $Y=26150
X372 1 M7_M6_CDNS_7651586358813 $T=74710 34150 0 0 $X=74350 $Y=34020
X373 1 M7_M6_CDNS_7651586358813 $T=74880 9920 0 0 $X=74520 $Y=9790
X374 2 M7_M6_CDNS_7651586358813 $T=77130 16720 0 0 $X=76770 $Y=16590
X375 2 M7_M6_CDNS_7651586358813 $T=77130 24150 0 0 $X=76770 $Y=24020
X376 2 M7_M6_CDNS_7651586358813 $T=77130 33380 0 0 $X=76770 $Y=33250
X377 2 M7_M6_CDNS_7651586358813 $T=78960 40520 0 0 $X=78600 $Y=40390
X378 1 M7_M6_CDNS_7651586358813 $T=83500 11170 0 0 $X=83140 $Y=11040
X379 1 M7_M6_CDNS_7651586358813 $T=85120 19020 0 0 $X=84760 $Y=18890
X380 1 M7_M6_CDNS_7651586358813 $T=85120 28370 0 0 $X=84760 $Y=28240
X381 1 M7_M6_CDNS_7651586358813 $T=85120 35150 0 0 $X=84760 $Y=35020
X382 2 M7_M6_CDNS_7651586358813 $T=99950 62120 0 0 $X=99590 $Y=61990
X383 2 M7_M6_CDNS_7651586358813 $T=100620 51980 0 0 $X=100260 $Y=51850
X384 2 M7_M6_CDNS_7651586358813 $T=102130 14020 0 0 $X=101770 $Y=13890
X385 2 M7_M6_CDNS_7651586358813 $T=102130 22060 0 0 $X=101770 $Y=21930
X386 2 M7_M6_CDNS_7651586358813 $T=102130 29250 0 0 $X=101770 $Y=29120
X387 2 M7_M6_CDNS_7651586358813 $T=102130 38320 0 0 $X=101770 $Y=38190
X388 2 M7_M6_CDNS_7651586358813 $T=105780 67340 0 0 $X=105420 $Y=67210
X389 1 M7_M6_CDNS_7651586358813 $T=106700 9920 0 0 $X=106340 $Y=9790
X390 1 M7_M6_CDNS_7651586358813 $T=106700 18310 0 0 $X=106340 $Y=18180
X391 1 M7_M6_CDNS_7651586358813 $T=106700 26700 0 0 $X=106340 $Y=26570
X392 1 M7_M6_CDNS_7651586358813 $T=106700 35090 0 0 $X=106340 $Y=34960
X393 1 M7_M6_CDNS_7651586358813 $T=106700 46070 0 0 $X=106340 $Y=45940
X394 1 M7_M6_CDNS_7651586358813 $T=106700 55950 0 0 $X=106340 $Y=55820
X395 1 M7_M6_CDNS_7651586358813 $T=106700 61400 0 0 $X=106340 $Y=61270
X396 1 M3_M2_CDNS_7651586358814 $T=17800 31900 0 0 $X=17440 $Y=31770
X397 1 M3_M2_CDNS_7651586358814 $T=17800 41260 0 0 $X=17440 $Y=41130
X398 1 M3_M2_CDNS_7651586358814 $T=17800 52820 0 0 $X=17440 $Y=52690
X399 1 M3_M2_CDNS_7651586358814 $T=17800 62680 0 0 $X=17440 $Y=62550
X400 2 M3_M2_CDNS_7651586358814 $T=19460 36430 0 0 $X=19100 $Y=36300
X401 2 M3_M2_CDNS_7651586358814 $T=19460 42880 0 0 $X=19100 $Y=42750
X402 2 M3_M2_CDNS_7651586358814 $T=19460 57580 0 0 $X=19100 $Y=57450
X403 2 M3_M2_CDNS_7651586358814 $T=19970 67840 0 0 $X=19610 $Y=67710
X404 1 M3_M2_CDNS_7651586358814 $T=25170 26030 0 0 $X=24810 $Y=25900
X405 1 M3_M2_CDNS_7651586358814 $T=25170 36370 0 0 $X=24810 $Y=36240
X406 1 M3_M2_CDNS_7651586358814 $T=26180 46210 0 0 $X=25820 $Y=46080
X407 1 M3_M2_CDNS_7651586358814 $T=26180 55960 0 0 $X=25820 $Y=55830
X408 2 M3_M2_CDNS_7651586358814 $T=29850 33170 0 0 $X=29490 $Y=33040
X409 2 M3_M2_CDNS_7651586358814 $T=29850 41710 0 0 $X=29490 $Y=41580
X410 2 M3_M2_CDNS_7651586358814 $T=29850 49920 0 0 $X=29490 $Y=49790
X411 2 M3_M2_CDNS_7651586358814 $T=29850 60150 0 0 $X=29490 $Y=60020
X412 1 M3_M2_CDNS_7651586358814 $T=31640 27290 0 0 $X=31280 $Y=27160
X413 1 M3_M2_CDNS_7651586358814 $T=31640 36130 0 0 $X=31280 $Y=36000
X414 1 M3_M2_CDNS_7651586358814 $T=31640 43470 0 0 $X=31280 $Y=43340
X415 1 M3_M2_CDNS_7651586358814 $T=31640 52000 0 0 $X=31280 $Y=51870
X416 1 M3_M2_CDNS_7651586358814 $T=47370 27010 0 0 $X=47010 $Y=26880
X417 1 M3_M2_CDNS_7651586358814 $T=47370 34360 0 0 $X=47010 $Y=34230
X418 1 M3_M2_CDNS_7651586358814 $T=48190 19140 0 0 $X=47830 $Y=19010
X419 1 M3_M2_CDNS_7651586358814 $T=50630 43060 0 0 $X=50270 $Y=42930
X420 2 M3_M2_CDNS_7651586358814 $T=52000 24420 0 0 $X=51640 $Y=24290
X421 2 M3_M2_CDNS_7651586358814 $T=52000 32940 0 0 $X=51640 $Y=32810
X422 2 M3_M2_CDNS_7651586358814 $T=52000 41710 0 0 $X=51640 $Y=41580
X423 2 M3_M2_CDNS_7651586358814 $T=52000 50750 0 0 $X=51640 $Y=50620
X424 2 M3_M2_CDNS_7651586358814 $T=52000 70000 0 0 $X=51640 $Y=69870
X425 1 M3_M2_CDNS_7651586358814 $T=54300 36130 0 0 $X=53940 $Y=36000
X426 1 M3_M2_CDNS_7651586358814 $T=57590 18970 0 0 $X=57230 $Y=18840
X427 1 M3_M2_CDNS_7651586358814 $T=57590 27180 0 0 $X=57230 $Y=27050
X428 1 M3_M2_CDNS_7651586358814 $T=58810 43370 0 0 $X=58450 $Y=43240
X429 1 M3_M2_CDNS_7651586358814 $T=74710 18350 0 0 $X=74350 $Y=18220
X430 1 M3_M2_CDNS_7651586358814 $T=74710 26280 0 0 $X=74350 $Y=26150
X431 1 M3_M2_CDNS_7651586358814 $T=74710 34150 0 0 $X=74350 $Y=34020
X432 1 M3_M2_CDNS_7651586358814 $T=74880 9920 0 0 $X=74520 $Y=9790
X433 2 M3_M2_CDNS_7651586358814 $T=77130 16720 0 0 $X=76770 $Y=16590
X434 2 M3_M2_CDNS_7651586358814 $T=77130 24150 0 0 $X=76770 $Y=24020
X435 2 M3_M2_CDNS_7651586358814 $T=77130 33380 0 0 $X=76770 $Y=33250
X436 2 M3_M2_CDNS_7651586358814 $T=78960 40520 0 0 $X=78600 $Y=40390
X437 1 M3_M2_CDNS_7651586358814 $T=83500 11170 0 0 $X=83140 $Y=11040
X438 1 M3_M2_CDNS_7651586358814 $T=85120 19020 0 0 $X=84760 $Y=18890
X439 1 M3_M2_CDNS_7651586358814 $T=85120 28370 0 0 $X=84760 $Y=28240
X440 1 M3_M2_CDNS_7651586358814 $T=85120 35150 0 0 $X=84760 $Y=35020
X441 2 M3_M2_CDNS_7651586358814 $T=99950 62120 0 0 $X=99590 $Y=61990
X442 2 M3_M2_CDNS_7651586358814 $T=100620 51980 0 0 $X=100260 $Y=51850
X443 2 M3_M2_CDNS_7651586358814 $T=102130 14020 0 0 $X=101770 $Y=13890
X444 2 M3_M2_CDNS_7651586358814 $T=102130 22060 0 0 $X=101770 $Y=21930
X445 2 M3_M2_CDNS_7651586358814 $T=102130 29250 0 0 $X=101770 $Y=29120
X446 2 M3_M2_CDNS_7651586358814 $T=102130 38320 0 0 $X=101770 $Y=38190
X447 2 M3_M2_CDNS_7651586358814 $T=105780 67340 0 0 $X=105420 $Y=67210
X448 1 M3_M2_CDNS_7651586358814 $T=106700 9920 0 0 $X=106340 $Y=9790
X449 1 M3_M2_CDNS_7651586358814 $T=106700 18310 0 0 $X=106340 $Y=18180
X450 1 M3_M2_CDNS_7651586358814 $T=106700 26700 0 0 $X=106340 $Y=26570
X451 1 M3_M2_CDNS_7651586358814 $T=106700 35090 0 0 $X=106340 $Y=34960
X452 1 M3_M2_CDNS_7651586358814 $T=106700 46070 0 0 $X=106340 $Y=45940
X453 1 M3_M2_CDNS_7651586358814 $T=106700 55950 0 0 $X=106340 $Y=55820
X454 1 M3_M2_CDNS_7651586358814 $T=106700 61400 0 0 $X=106340 $Y=61270
X455 46 M3_M2_CDNS_7651586358815 $T=83660 14830 0 0 $X=83440 $Y=14700
X456 46 M3_M2_CDNS_7651586358815 $T=83660 22300 0 0 $X=83440 $Y=22170
X457 46 M3_M2_CDNS_7651586358815 $T=83660 31480 0 0 $X=83440 $Y=31350
X458 46 M3_M2_CDNS_7651586358815 $T=83660 38710 0 0 $X=83440 $Y=38580
X459 47 M3_M2_CDNS_7651586358815 $T=91230 14480 0 0 $X=91010 $Y=14350
X460 47 M3_M2_CDNS_7651586358815 $T=91230 21950 0 0 $X=91010 $Y=21820
X461 47 M3_M2_CDNS_7651586358815 $T=91230 31130 0 0 $X=91010 $Y=31000
X462 47 M3_M2_CDNS_7651586358815 $T=91230 38320 0 0 $X=91010 $Y=38190
X463 48 M3_M2_CDNS_7651586358815 $T=92110 15580 0 0 $X=91890 $Y=15450
X464 49 M3_M2_CDNS_7651586358815 $T=92110 23050 0 0 $X=91890 $Y=22920
X465 50 M3_M2_CDNS_7651586358815 $T=92110 32230 0 0 $X=91890 $Y=32100
X466 51 M3_M2_CDNS_7651586358815 $T=92110 39460 0 0 $X=91890 $Y=39330
X467 46 M3_M2_CDNS_7651586358815 $T=93260 10940 0 0 $X=93040 $Y=10810
X468 46 M3_M2_CDNS_7651586358815 $T=93260 18410 0 0 $X=93040 $Y=18280
X469 46 M3_M2_CDNS_7651586358815 $T=93260 27590 0 0 $X=93040 $Y=27460
X470 46 M3_M2_CDNS_7651586358815 $T=93260 34820 0 0 $X=93040 $Y=34690
X471 46 M3_M2_CDNS_7651586358815 $T=99520 48720 0 0 $X=99300 $Y=48590
X472 46 M3_M2_CDNS_7651586358815 $T=99520 58720 0 0 $X=99300 $Y=58590
X473 47 M3_M2_CDNS_7651586358815 $T=100830 10590 0 0 $X=100610 $Y=10460
X474 47 M3_M2_CDNS_7651586358815 $T=100830 18060 0 0 $X=100610 $Y=17930
X475 47 M3_M2_CDNS_7651586358815 $T=100830 27240 0 0 $X=100610 $Y=27110
X476 47 M3_M2_CDNS_7651586358815 $T=100830 34470 0 0 $X=100610 $Y=34340
X477 52 M3_M2_CDNS_7651586358815 $T=101710 11690 0 0 $X=101490 $Y=11560
X478 53 M3_M2_CDNS_7651586358815 $T=101710 19160 0 0 $X=101490 $Y=19030
X479 54 M3_M2_CDNS_7651586358815 $T=101710 28340 0 0 $X=101490 $Y=28210
X480 55 M3_M2_CDNS_7651586358815 $T=101710 35570 0 0 $X=101490 $Y=35440
X481 46 M3_M2_CDNS_7651586358815 $T=104930 64130 0 0 $X=104710 $Y=64000
X482 47 M3_M2_CDNS_7651586358815 $T=107050 58360 0 0 $X=106830 $Y=58230
X483 47 M3_M2_CDNS_7651586358815 $T=107080 48320 0 0 $X=106860 $Y=48190
X484 56 M3_M2_CDNS_7651586358815 $T=107970 49470 0 0 $X=107750 $Y=49340
X485 57 M3_M2_CDNS_7651586358815 $T=107970 59470 0 0 $X=107750 $Y=59340
X486 47 M3_M2_CDNS_7651586358815 $T=112490 63750 0 0 $X=112270 $Y=63620
X487 58 M3_M2_CDNS_7651586358815 $T=113380 64880 0 0 $X=113160 $Y=64750
X488 1 M8_M7_CDNS_7651586358816 $T=17800 31900 0 0 $X=17440 $Y=31770
X489 1 M8_M7_CDNS_7651586358816 $T=17800 41260 0 0 $X=17440 $Y=41130
X490 1 M8_M7_CDNS_7651586358816 $T=17800 52820 0 0 $X=17440 $Y=52690
X491 1 M8_M7_CDNS_7651586358816 $T=17800 62680 0 0 $X=17440 $Y=62550
X492 2 M8_M7_CDNS_7651586358816 $T=19460 36430 0 0 $X=19100 $Y=36300
X493 2 M8_M7_CDNS_7651586358816 $T=19460 42880 0 0 $X=19100 $Y=42750
X494 2 M8_M7_CDNS_7651586358816 $T=19460 57580 0 0 $X=19100 $Y=57450
X495 2 M8_M7_CDNS_7651586358816 $T=19970 67840 0 0 $X=19610 $Y=67710
X496 1 M8_M7_CDNS_7651586358816 $T=25170 26030 0 0 $X=24810 $Y=25900
X497 1 M8_M7_CDNS_7651586358816 $T=25170 36370 0 0 $X=24810 $Y=36240
X498 1 M8_M7_CDNS_7651586358816 $T=26180 46210 0 0 $X=25820 $Y=46080
X499 1 M8_M7_CDNS_7651586358816 $T=26180 55960 0 0 $X=25820 $Y=55830
X500 2 M8_M7_CDNS_7651586358816 $T=29850 33170 0 0 $X=29490 $Y=33040
X501 2 M8_M7_CDNS_7651586358816 $T=29850 41710 0 0 $X=29490 $Y=41580
X502 2 M8_M7_CDNS_7651586358816 $T=29850 49920 0 0 $X=29490 $Y=49790
X503 2 M8_M7_CDNS_7651586358816 $T=29850 60150 0 0 $X=29490 $Y=60020
X504 1 M8_M7_CDNS_7651586358816 $T=31640 27290 0 0 $X=31280 $Y=27160
X505 1 M8_M7_CDNS_7651586358816 $T=31640 36130 0 0 $X=31280 $Y=36000
X506 1 M8_M7_CDNS_7651586358816 $T=31640 43470 0 0 $X=31280 $Y=43340
X507 1 M8_M7_CDNS_7651586358816 $T=31640 52000 0 0 $X=31280 $Y=51870
X508 1 M8_M7_CDNS_7651586358816 $T=47370 27010 0 0 $X=47010 $Y=26880
X509 1 M8_M7_CDNS_7651586358816 $T=47370 34360 0 0 $X=47010 $Y=34230
X510 1 M8_M7_CDNS_7651586358816 $T=48190 19140 0 0 $X=47830 $Y=19010
X511 1 M8_M7_CDNS_7651586358816 $T=50630 43060 0 0 $X=50270 $Y=42930
X512 2 M8_M7_CDNS_7651586358816 $T=52000 24420 0 0 $X=51640 $Y=24290
X513 2 M8_M7_CDNS_7651586358816 $T=52000 32940 0 0 $X=51640 $Y=32810
X514 2 M8_M7_CDNS_7651586358816 $T=52000 41710 0 0 $X=51640 $Y=41580
X515 2 M8_M7_CDNS_7651586358816 $T=52000 50750 0 0 $X=51640 $Y=50620
X516 2 M8_M7_CDNS_7651586358816 $T=52000 70000 0 0 $X=51640 $Y=69870
X517 1 M8_M7_CDNS_7651586358816 $T=54300 36130 0 0 $X=53940 $Y=36000
X518 1 M8_M7_CDNS_7651586358816 $T=57590 18970 0 0 $X=57230 $Y=18840
X519 1 M8_M7_CDNS_7651586358816 $T=57590 27180 0 0 $X=57230 $Y=27050
X520 1 M8_M7_CDNS_7651586358816 $T=58810 43370 0 0 $X=58450 $Y=43240
X521 1 M8_M7_CDNS_7651586358816 $T=74710 18350 0 0 $X=74350 $Y=18220
X522 1 M8_M7_CDNS_7651586358816 $T=74710 26280 0 0 $X=74350 $Y=26150
X523 1 M8_M7_CDNS_7651586358816 $T=74710 34150 0 0 $X=74350 $Y=34020
X524 1 M8_M7_CDNS_7651586358816 $T=74880 9920 0 0 $X=74520 $Y=9790
X525 2 M8_M7_CDNS_7651586358816 $T=77130 16720 0 0 $X=76770 $Y=16590
X526 2 M8_M7_CDNS_7651586358816 $T=77130 24150 0 0 $X=76770 $Y=24020
X527 2 M8_M7_CDNS_7651586358816 $T=77130 33380 0 0 $X=76770 $Y=33250
X528 2 M8_M7_CDNS_7651586358816 $T=78960 40520 0 0 $X=78600 $Y=40390
X529 1 M8_M7_CDNS_7651586358816 $T=83500 11170 0 0 $X=83140 $Y=11040
X530 1 M8_M7_CDNS_7651586358816 $T=85120 19020 0 0 $X=84760 $Y=18890
X531 1 M8_M7_CDNS_7651586358816 $T=85120 28370 0 0 $X=84760 $Y=28240
X532 1 M8_M7_CDNS_7651586358816 $T=85120 35150 0 0 $X=84760 $Y=35020
X533 2 M8_M7_CDNS_7651586358816 $T=99950 62120 0 0 $X=99590 $Y=61990
X534 2 M8_M7_CDNS_7651586358816 $T=100620 51980 0 0 $X=100260 $Y=51850
X535 2 M8_M7_CDNS_7651586358816 $T=102130 14020 0 0 $X=101770 $Y=13890
X536 2 M8_M7_CDNS_7651586358816 $T=102130 22060 0 0 $X=101770 $Y=21930
X537 2 M8_M7_CDNS_7651586358816 $T=102130 29250 0 0 $X=101770 $Y=29120
X538 2 M8_M7_CDNS_7651586358816 $T=102130 38320 0 0 $X=101770 $Y=38190
X539 2 M8_M7_CDNS_7651586358816 $T=105780 67340 0 0 $X=105420 $Y=67210
X540 1 M8_M7_CDNS_7651586358816 $T=106700 9920 0 0 $X=106340 $Y=9790
X541 1 M8_M7_CDNS_7651586358816 $T=106700 18310 0 0 $X=106340 $Y=18180
X542 1 M8_M7_CDNS_7651586358816 $T=106700 26700 0 0 $X=106340 $Y=26570
X543 1 M8_M7_CDNS_7651586358816 $T=106700 35090 0 0 $X=106340 $Y=34960
X544 1 M8_M7_CDNS_7651586358816 $T=106700 46070 0 0 $X=106340 $Y=45940
X545 1 M8_M7_CDNS_7651586358816 $T=106700 55950 0 0 $X=106340 $Y=55820
X546 1 M8_M7_CDNS_7651586358816 $T=106700 61400 0 0 $X=106340 $Y=61270
X547 1 M2_M1_CDNS_7651586358817 $T=17800 31900 0 0 $X=17440 $Y=31770
X548 1 M2_M1_CDNS_7651586358817 $T=17800 41260 0 0 $X=17440 $Y=41130
X549 1 M2_M1_CDNS_7651586358817 $T=17800 52820 0 0 $X=17440 $Y=52690
X550 1 M2_M1_CDNS_7651586358817 $T=17800 62680 0 0 $X=17440 $Y=62550
X551 2 M2_M1_CDNS_7651586358817 $T=19460 36430 0 0 $X=19100 $Y=36300
X552 2 M2_M1_CDNS_7651586358817 $T=19460 42880 0 0 $X=19100 $Y=42750
X553 2 M2_M1_CDNS_7651586358817 $T=19460 57580 0 0 $X=19100 $Y=57450
X554 2 M2_M1_CDNS_7651586358817 $T=19970 67840 0 0 $X=19610 $Y=67710
X555 1 M2_M1_CDNS_7651586358817 $T=25170 26030 0 0 $X=24810 $Y=25900
X556 1 M2_M1_CDNS_7651586358817 $T=25170 36370 0 0 $X=24810 $Y=36240
X557 1 M2_M1_CDNS_7651586358817 $T=26180 46210 0 0 $X=25820 $Y=46080
X558 1 M2_M1_CDNS_7651586358817 $T=26180 55960 0 0 $X=25820 $Y=55830
X559 2 M2_M1_CDNS_7651586358817 $T=29850 33170 0 0 $X=29490 $Y=33040
X560 2 M2_M1_CDNS_7651586358817 $T=29850 41710 0 0 $X=29490 $Y=41580
X561 2 M2_M1_CDNS_7651586358817 $T=29850 49920 0 0 $X=29490 $Y=49790
X562 2 M2_M1_CDNS_7651586358817 $T=29850 60150 0 0 $X=29490 $Y=60020
X563 1 M2_M1_CDNS_7651586358817 $T=31640 27290 0 0 $X=31280 $Y=27160
X564 1 M2_M1_CDNS_7651586358817 $T=31640 36130 0 0 $X=31280 $Y=36000
X565 1 M2_M1_CDNS_7651586358817 $T=31640 43470 0 0 $X=31280 $Y=43340
X566 1 M2_M1_CDNS_7651586358817 $T=31640 52000 0 0 $X=31280 $Y=51870
X567 1 M2_M1_CDNS_7651586358817 $T=47370 27010 0 0 $X=47010 $Y=26880
X568 1 M2_M1_CDNS_7651586358817 $T=47370 34360 0 0 $X=47010 $Y=34230
X569 1 M2_M1_CDNS_7651586358817 $T=48190 19140 0 0 $X=47830 $Y=19010
X570 1 M2_M1_CDNS_7651586358817 $T=50630 43060 0 0 $X=50270 $Y=42930
X571 2 M2_M1_CDNS_7651586358817 $T=52000 24420 0 0 $X=51640 $Y=24290
X572 2 M2_M1_CDNS_7651586358817 $T=52000 32940 0 0 $X=51640 $Y=32810
X573 2 M2_M1_CDNS_7651586358817 $T=52000 41710 0 0 $X=51640 $Y=41580
X574 2 M2_M1_CDNS_7651586358817 $T=52000 50750 0 0 $X=51640 $Y=50620
X575 2 M2_M1_CDNS_7651586358817 $T=52000 70000 0 0 $X=51640 $Y=69870
X576 1 M2_M1_CDNS_7651586358817 $T=54300 36130 0 0 $X=53940 $Y=36000
X577 1 M2_M1_CDNS_7651586358817 $T=57590 18970 0 0 $X=57230 $Y=18840
X578 1 M2_M1_CDNS_7651586358817 $T=57590 27180 0 0 $X=57230 $Y=27050
X579 1 M2_M1_CDNS_7651586358817 $T=58810 43370 0 0 $X=58450 $Y=43240
X580 1 M2_M1_CDNS_7651586358817 $T=74710 18350 0 0 $X=74350 $Y=18220
X581 1 M2_M1_CDNS_7651586358817 $T=74710 26280 0 0 $X=74350 $Y=26150
X582 1 M2_M1_CDNS_7651586358817 $T=74710 34150 0 0 $X=74350 $Y=34020
X583 1 M2_M1_CDNS_7651586358817 $T=74880 9920 0 0 $X=74520 $Y=9790
X584 2 M2_M1_CDNS_7651586358817 $T=77130 16720 0 0 $X=76770 $Y=16590
X585 2 M2_M1_CDNS_7651586358817 $T=77130 24150 0 0 $X=76770 $Y=24020
X586 2 M2_M1_CDNS_7651586358817 $T=77130 33380 0 0 $X=76770 $Y=33250
X587 2 M2_M1_CDNS_7651586358817 $T=78960 40520 0 0 $X=78600 $Y=40390
X588 1 M2_M1_CDNS_7651586358817 $T=83500 11170 0 0 $X=83140 $Y=11040
X589 1 M2_M1_CDNS_7651586358817 $T=85120 19020 0 0 $X=84760 $Y=18890
X590 1 M2_M1_CDNS_7651586358817 $T=85120 28370 0 0 $X=84760 $Y=28240
X591 1 M2_M1_CDNS_7651586358817 $T=85120 35150 0 0 $X=84760 $Y=35020
X592 2 M2_M1_CDNS_7651586358817 $T=99950 62120 0 0 $X=99590 $Y=61990
X593 2 M2_M1_CDNS_7651586358817 $T=100620 51980 0 0 $X=100260 $Y=51850
X594 2 M2_M1_CDNS_7651586358817 $T=102130 14020 0 0 $X=101770 $Y=13890
X595 2 M2_M1_CDNS_7651586358817 $T=102130 22060 0 0 $X=101770 $Y=21930
X596 2 M2_M1_CDNS_7651586358817 $T=102130 29250 0 0 $X=101770 $Y=29120
X597 2 M2_M1_CDNS_7651586358817 $T=102130 38320 0 0 $X=101770 $Y=38190
X598 2 M2_M1_CDNS_7651586358817 $T=105780 67340 0 0 $X=105420 $Y=67210
X599 1 M2_M1_CDNS_7651586358817 $T=106700 9920 0 0 $X=106340 $Y=9790
X600 1 M2_M1_CDNS_7651586358817 $T=106700 18310 0 0 $X=106340 $Y=18180
X601 1 M2_M1_CDNS_7651586358817 $T=106700 26700 0 0 $X=106340 $Y=26570
X602 1 M2_M1_CDNS_7651586358817 $T=106700 35090 0 0 $X=106340 $Y=34960
X603 1 M2_M1_CDNS_7651586358817 $T=106700 46070 0 0 $X=106340 $Y=45940
X604 1 M2_M1_CDNS_7651586358817 $T=106700 55950 0 0 $X=106340 $Y=55820
X605 1 M2_M1_CDNS_7651586358817 $T=106700 61400 0 0 $X=106340 $Y=61270
X606 1 M4_M3_CDNS_7651586358818 $T=17800 31900 0 0 $X=17440 $Y=31770
X607 1 M4_M3_CDNS_7651586358818 $T=17800 41260 0 0 $X=17440 $Y=41130
X608 1 M4_M3_CDNS_7651586358818 $T=17800 52820 0 0 $X=17440 $Y=52690
X609 1 M4_M3_CDNS_7651586358818 $T=17800 62680 0 0 $X=17440 $Y=62550
X610 2 M4_M3_CDNS_7651586358818 $T=19460 36430 0 0 $X=19100 $Y=36300
X611 2 M4_M3_CDNS_7651586358818 $T=19460 42880 0 0 $X=19100 $Y=42750
X612 2 M4_M3_CDNS_7651586358818 $T=19460 57580 0 0 $X=19100 $Y=57450
X613 2 M4_M3_CDNS_7651586358818 $T=19970 67840 0 0 $X=19610 $Y=67710
X614 1 M4_M3_CDNS_7651586358818 $T=25170 26030 0 0 $X=24810 $Y=25900
X615 1 M4_M3_CDNS_7651586358818 $T=25170 36370 0 0 $X=24810 $Y=36240
X616 1 M4_M3_CDNS_7651586358818 $T=26180 46210 0 0 $X=25820 $Y=46080
X617 1 M4_M3_CDNS_7651586358818 $T=26180 55960 0 0 $X=25820 $Y=55830
X618 2 M4_M3_CDNS_7651586358818 $T=29850 33170 0 0 $X=29490 $Y=33040
X619 2 M4_M3_CDNS_7651586358818 $T=29850 41710 0 0 $X=29490 $Y=41580
X620 2 M4_M3_CDNS_7651586358818 $T=29850 49920 0 0 $X=29490 $Y=49790
X621 2 M4_M3_CDNS_7651586358818 $T=29850 60150 0 0 $X=29490 $Y=60020
X622 1 M4_M3_CDNS_7651586358818 $T=31640 27290 0 0 $X=31280 $Y=27160
X623 1 M4_M3_CDNS_7651586358818 $T=31640 36130 0 0 $X=31280 $Y=36000
X624 1 M4_M3_CDNS_7651586358818 $T=31640 43470 0 0 $X=31280 $Y=43340
X625 1 M4_M3_CDNS_7651586358818 $T=31640 52000 0 0 $X=31280 $Y=51870
X626 1 M4_M3_CDNS_7651586358818 $T=47370 27010 0 0 $X=47010 $Y=26880
X627 1 M4_M3_CDNS_7651586358818 $T=47370 34360 0 0 $X=47010 $Y=34230
X628 1 M4_M3_CDNS_7651586358818 $T=48190 19140 0 0 $X=47830 $Y=19010
X629 1 M4_M3_CDNS_7651586358818 $T=50630 43060 0 0 $X=50270 $Y=42930
X630 2 M4_M3_CDNS_7651586358818 $T=52000 24420 0 0 $X=51640 $Y=24290
X631 2 M4_M3_CDNS_7651586358818 $T=52000 32940 0 0 $X=51640 $Y=32810
X632 2 M4_M3_CDNS_7651586358818 $T=52000 41710 0 0 $X=51640 $Y=41580
X633 2 M4_M3_CDNS_7651586358818 $T=52000 50750 0 0 $X=51640 $Y=50620
X634 2 M4_M3_CDNS_7651586358818 $T=52000 70000 0 0 $X=51640 $Y=69870
X635 1 M4_M3_CDNS_7651586358818 $T=54300 36130 0 0 $X=53940 $Y=36000
X636 1 M4_M3_CDNS_7651586358818 $T=57590 18970 0 0 $X=57230 $Y=18840
X637 1 M4_M3_CDNS_7651586358818 $T=57590 27180 0 0 $X=57230 $Y=27050
X638 1 M4_M3_CDNS_7651586358818 $T=58810 43370 0 0 $X=58450 $Y=43240
X639 1 M4_M3_CDNS_7651586358818 $T=74710 18350 0 0 $X=74350 $Y=18220
X640 1 M4_M3_CDNS_7651586358818 $T=74710 26280 0 0 $X=74350 $Y=26150
X641 1 M4_M3_CDNS_7651586358818 $T=74710 34150 0 0 $X=74350 $Y=34020
X642 1 M4_M3_CDNS_7651586358818 $T=74880 9920 0 0 $X=74520 $Y=9790
X643 2 M4_M3_CDNS_7651586358818 $T=77130 16720 0 0 $X=76770 $Y=16590
X644 2 M4_M3_CDNS_7651586358818 $T=77130 24150 0 0 $X=76770 $Y=24020
X645 2 M4_M3_CDNS_7651586358818 $T=77130 33380 0 0 $X=76770 $Y=33250
X646 2 M4_M3_CDNS_7651586358818 $T=78960 40520 0 0 $X=78600 $Y=40390
X647 1 M4_M3_CDNS_7651586358818 $T=83500 11170 0 0 $X=83140 $Y=11040
X648 1 M4_M3_CDNS_7651586358818 $T=85120 19020 0 0 $X=84760 $Y=18890
X649 1 M4_M3_CDNS_7651586358818 $T=85120 28370 0 0 $X=84760 $Y=28240
X650 1 M4_M3_CDNS_7651586358818 $T=85120 35150 0 0 $X=84760 $Y=35020
X651 2 M4_M3_CDNS_7651586358818 $T=99950 62120 0 0 $X=99590 $Y=61990
X652 2 M4_M3_CDNS_7651586358818 $T=100620 51980 0 0 $X=100260 $Y=51850
X653 2 M4_M3_CDNS_7651586358818 $T=102130 14020 0 0 $X=101770 $Y=13890
X654 2 M4_M3_CDNS_7651586358818 $T=102130 22060 0 0 $X=101770 $Y=21930
X655 2 M4_M3_CDNS_7651586358818 $T=102130 29250 0 0 $X=101770 $Y=29120
X656 2 M4_M3_CDNS_7651586358818 $T=102130 38320 0 0 $X=101770 $Y=38190
X657 2 M4_M3_CDNS_7651586358818 $T=105780 67340 0 0 $X=105420 $Y=67210
X658 1 M4_M3_CDNS_7651586358818 $T=106700 9920 0 0 $X=106340 $Y=9790
X659 1 M4_M3_CDNS_7651586358818 $T=106700 18310 0 0 $X=106340 $Y=18180
X660 1 M4_M3_CDNS_7651586358818 $T=106700 26700 0 0 $X=106340 $Y=26570
X661 1 M4_M3_CDNS_7651586358818 $T=106700 35090 0 0 $X=106340 $Y=34960
X662 1 M4_M3_CDNS_7651586358818 $T=106700 46070 0 0 $X=106340 $Y=45940
X663 1 M4_M3_CDNS_7651586358818 $T=106700 55950 0 0 $X=106340 $Y=55820
X664 1 M4_M3_CDNS_7651586358818 $T=106700 61400 0 0 $X=106340 $Y=61270
X665 1 M6_M5_CDNS_7651586358819 $T=17800 31900 0 0 $X=17440 $Y=31770
X666 1 M6_M5_CDNS_7651586358819 $T=17800 41260 0 0 $X=17440 $Y=41130
X667 1 M6_M5_CDNS_7651586358819 $T=17800 52820 0 0 $X=17440 $Y=52690
X668 1 M6_M5_CDNS_7651586358819 $T=17800 62680 0 0 $X=17440 $Y=62550
X669 2 M6_M5_CDNS_7651586358819 $T=19460 36430 0 0 $X=19100 $Y=36300
X670 2 M6_M5_CDNS_7651586358819 $T=19460 42880 0 0 $X=19100 $Y=42750
X671 2 M6_M5_CDNS_7651586358819 $T=19460 57580 0 0 $X=19100 $Y=57450
X672 2 M6_M5_CDNS_7651586358819 $T=19970 67840 0 0 $X=19610 $Y=67710
X673 1 M6_M5_CDNS_7651586358819 $T=25170 26030 0 0 $X=24810 $Y=25900
X674 1 M6_M5_CDNS_7651586358819 $T=25170 36370 0 0 $X=24810 $Y=36240
X675 1 M6_M5_CDNS_7651586358819 $T=26180 46210 0 0 $X=25820 $Y=46080
X676 1 M6_M5_CDNS_7651586358819 $T=26180 55960 0 0 $X=25820 $Y=55830
X677 2 M6_M5_CDNS_7651586358819 $T=29850 33170 0 0 $X=29490 $Y=33040
X678 2 M6_M5_CDNS_7651586358819 $T=29850 41710 0 0 $X=29490 $Y=41580
X679 2 M6_M5_CDNS_7651586358819 $T=29850 49920 0 0 $X=29490 $Y=49790
X680 2 M6_M5_CDNS_7651586358819 $T=29850 60150 0 0 $X=29490 $Y=60020
X681 1 M6_M5_CDNS_7651586358819 $T=31640 27290 0 0 $X=31280 $Y=27160
X682 1 M6_M5_CDNS_7651586358819 $T=31640 36130 0 0 $X=31280 $Y=36000
X683 1 M6_M5_CDNS_7651586358819 $T=31640 43470 0 0 $X=31280 $Y=43340
X684 1 M6_M5_CDNS_7651586358819 $T=31640 52000 0 0 $X=31280 $Y=51870
X685 1 M6_M5_CDNS_7651586358819 $T=47370 27010 0 0 $X=47010 $Y=26880
X686 1 M6_M5_CDNS_7651586358819 $T=47370 34360 0 0 $X=47010 $Y=34230
X687 1 M6_M5_CDNS_7651586358819 $T=48190 19140 0 0 $X=47830 $Y=19010
X688 1 M6_M5_CDNS_7651586358819 $T=50630 43060 0 0 $X=50270 $Y=42930
X689 2 M6_M5_CDNS_7651586358819 $T=52000 24420 0 0 $X=51640 $Y=24290
X690 2 M6_M5_CDNS_7651586358819 $T=52000 32940 0 0 $X=51640 $Y=32810
X691 2 M6_M5_CDNS_7651586358819 $T=52000 41710 0 0 $X=51640 $Y=41580
X692 2 M6_M5_CDNS_7651586358819 $T=52000 50750 0 0 $X=51640 $Y=50620
X693 2 M6_M5_CDNS_7651586358819 $T=52000 70000 0 0 $X=51640 $Y=69870
X694 1 M6_M5_CDNS_7651586358819 $T=54300 36130 0 0 $X=53940 $Y=36000
X695 1 M6_M5_CDNS_7651586358819 $T=57590 18970 0 0 $X=57230 $Y=18840
X696 1 M6_M5_CDNS_7651586358819 $T=57590 27180 0 0 $X=57230 $Y=27050
X697 1 M6_M5_CDNS_7651586358819 $T=58810 43370 0 0 $X=58450 $Y=43240
X698 1 M6_M5_CDNS_7651586358819 $T=74710 18350 0 0 $X=74350 $Y=18220
X699 1 M6_M5_CDNS_7651586358819 $T=74710 26280 0 0 $X=74350 $Y=26150
X700 1 M6_M5_CDNS_7651586358819 $T=74710 34150 0 0 $X=74350 $Y=34020
X701 1 M6_M5_CDNS_7651586358819 $T=74880 9920 0 0 $X=74520 $Y=9790
X702 2 M6_M5_CDNS_7651586358819 $T=77130 16720 0 0 $X=76770 $Y=16590
X703 2 M6_M5_CDNS_7651586358819 $T=77130 24150 0 0 $X=76770 $Y=24020
X704 2 M6_M5_CDNS_7651586358819 $T=77130 33380 0 0 $X=76770 $Y=33250
X705 2 M6_M5_CDNS_7651586358819 $T=78960 40520 0 0 $X=78600 $Y=40390
X706 1 M6_M5_CDNS_7651586358819 $T=83500 11170 0 0 $X=83140 $Y=11040
X707 1 M6_M5_CDNS_7651586358819 $T=85120 19020 0 0 $X=84760 $Y=18890
X708 1 M6_M5_CDNS_7651586358819 $T=85120 28370 0 0 $X=84760 $Y=28240
X709 1 M6_M5_CDNS_7651586358819 $T=85120 35150 0 0 $X=84760 $Y=35020
X710 2 M6_M5_CDNS_7651586358819 $T=99950 62120 0 0 $X=99590 $Y=61990
X711 2 M6_M5_CDNS_7651586358819 $T=100620 51980 0 0 $X=100260 $Y=51850
X712 2 M6_M5_CDNS_7651586358819 $T=102130 14020 0 0 $X=101770 $Y=13890
X713 2 M6_M5_CDNS_7651586358819 $T=102130 22060 0 0 $X=101770 $Y=21930
X714 2 M6_M5_CDNS_7651586358819 $T=102130 29250 0 0 $X=101770 $Y=29120
X715 2 M6_M5_CDNS_7651586358819 $T=102130 38320 0 0 $X=101770 $Y=38190
X716 2 M6_M5_CDNS_7651586358819 $T=105780 67340 0 0 $X=105420 $Y=67210
X717 1 M6_M5_CDNS_7651586358819 $T=106700 9920 0 0 $X=106340 $Y=9790
X718 1 M6_M5_CDNS_7651586358819 $T=106700 18310 0 0 $X=106340 $Y=18180
X719 1 M6_M5_CDNS_7651586358819 $T=106700 26700 0 0 $X=106340 $Y=26570
X720 1 M6_M5_CDNS_7651586358819 $T=106700 35090 0 0 $X=106340 $Y=34960
X721 1 M6_M5_CDNS_7651586358819 $T=106700 46070 0 0 $X=106340 $Y=45940
X722 1 M6_M5_CDNS_7651586358819 $T=106700 55950 0 0 $X=106340 $Y=55820
X723 1 M6_M5_CDNS_7651586358819 $T=106700 61400 0 0 $X=106340 $Y=61270
X724 47 M2_M1_CDNS_7651586358820 $T=91230 14480 0 0 $X=91010 $Y=14350
X725 47 M2_M1_CDNS_7651586358820 $T=91230 21950 0 0 $X=91010 $Y=21820
X726 47 M2_M1_CDNS_7651586358820 $T=91230 31130 0 0 $X=91010 $Y=31000
X727 47 M2_M1_CDNS_7651586358820 $T=91230 38320 0 0 $X=91010 $Y=38190
X728 48 M2_M1_CDNS_7651586358820 $T=92110 15580 0 0 $X=91890 $Y=15450
X729 49 M2_M1_CDNS_7651586358820 $T=92110 23050 0 0 $X=91890 $Y=22920
X730 50 M2_M1_CDNS_7651586358820 $T=92110 32230 0 0 $X=91890 $Y=32100
X731 51 M2_M1_CDNS_7651586358820 $T=92110 39460 0 0 $X=91890 $Y=39330
X732 47 M2_M1_CDNS_7651586358820 $T=100830 10590 0 0 $X=100610 $Y=10460
X733 47 M2_M1_CDNS_7651586358820 $T=100830 18060 0 0 $X=100610 $Y=17930
X734 47 M2_M1_CDNS_7651586358820 $T=100830 27240 0 0 $X=100610 $Y=27110
X735 47 M2_M1_CDNS_7651586358820 $T=100830 34470 0 0 $X=100610 $Y=34340
X736 52 M2_M1_CDNS_7651586358820 $T=101710 11690 0 0 $X=101490 $Y=11560
X737 53 M2_M1_CDNS_7651586358820 $T=101710 19160 0 0 $X=101490 $Y=19030
X738 54 M2_M1_CDNS_7651586358820 $T=101710 28340 0 0 $X=101490 $Y=28210
X739 55 M2_M1_CDNS_7651586358820 $T=101710 35570 0 0 $X=101490 $Y=35440
X740 47 M2_M1_CDNS_7651586358820 $T=107050 58360 0 0 $X=106830 $Y=58230
X741 47 M2_M1_CDNS_7651586358820 $T=107080 48320 0 0 $X=106860 $Y=48190
X742 56 M2_M1_CDNS_7651586358820 $T=107970 49470 0 0 $X=107750 $Y=49340
X743 57 M2_M1_CDNS_7651586358820 $T=107970 59470 0 0 $X=107750 $Y=59340
X744 47 M2_M1_CDNS_7651586358820 $T=112490 63750 0 0 $X=112270 $Y=63620
X745 58 M2_M1_CDNS_7651586358820 $T=113380 64880 0 0 $X=113160 $Y=64750
X746 1 M9_M8_CDNS_7651586358821 $T=17800 31900 0 0 $X=17440 $Y=31770
X747 1 M9_M8_CDNS_7651586358821 $T=17800 41260 0 0 $X=17440 $Y=41130
X748 1 M9_M8_CDNS_7651586358821 $T=17800 52820 0 0 $X=17440 $Y=52690
X749 1 M9_M8_CDNS_7651586358821 $T=17800 62680 0 0 $X=17440 $Y=62550
X750 2 M9_M8_CDNS_7651586358821 $T=19460 36430 0 0 $X=19100 $Y=36300
X751 2 M9_M8_CDNS_7651586358821 $T=19460 42880 0 0 $X=19100 $Y=42750
X752 2 M9_M8_CDNS_7651586358821 $T=19460 57580 0 0 $X=19100 $Y=57450
X753 2 M9_M8_CDNS_7651586358821 $T=19970 67840 0 0 $X=19610 $Y=67710
X754 1 M9_M8_CDNS_7651586358821 $T=25170 26030 0 0 $X=24810 $Y=25900
X755 1 M9_M8_CDNS_7651586358821 $T=25170 36370 0 0 $X=24810 $Y=36240
X756 1 M9_M8_CDNS_7651586358821 $T=26180 46210 0 0 $X=25820 $Y=46080
X757 1 M9_M8_CDNS_7651586358821 $T=26180 55960 0 0 $X=25820 $Y=55830
X758 2 M9_M8_CDNS_7651586358821 $T=29850 33170 0 0 $X=29490 $Y=33040
X759 2 M9_M8_CDNS_7651586358821 $T=29850 41710 0 0 $X=29490 $Y=41580
X760 2 M9_M8_CDNS_7651586358821 $T=29850 49920 0 0 $X=29490 $Y=49790
X761 2 M9_M8_CDNS_7651586358821 $T=29850 60150 0 0 $X=29490 $Y=60020
X762 1 M9_M8_CDNS_7651586358821 $T=31640 27290 0 0 $X=31280 $Y=27160
X763 1 M9_M8_CDNS_7651586358821 $T=31640 36130 0 0 $X=31280 $Y=36000
X764 1 M9_M8_CDNS_7651586358821 $T=31640 43470 0 0 $X=31280 $Y=43340
X765 1 M9_M8_CDNS_7651586358821 $T=31640 52000 0 0 $X=31280 $Y=51870
X766 1 M9_M8_CDNS_7651586358821 $T=47370 27010 0 0 $X=47010 $Y=26880
X767 1 M9_M8_CDNS_7651586358821 $T=47370 34360 0 0 $X=47010 $Y=34230
X768 1 M9_M8_CDNS_7651586358821 $T=48190 19140 0 0 $X=47830 $Y=19010
X769 1 M9_M8_CDNS_7651586358821 $T=50630 43060 0 0 $X=50270 $Y=42930
X770 2 M9_M8_CDNS_7651586358821 $T=52000 24420 0 0 $X=51640 $Y=24290
X771 2 M9_M8_CDNS_7651586358821 $T=52000 32940 0 0 $X=51640 $Y=32810
X772 2 M9_M8_CDNS_7651586358821 $T=52000 41710 0 0 $X=51640 $Y=41580
X773 2 M9_M8_CDNS_7651586358821 $T=52000 50750 0 0 $X=51640 $Y=50620
X774 2 M9_M8_CDNS_7651586358821 $T=52000 70000 0 0 $X=51640 $Y=69870
X775 1 M9_M8_CDNS_7651586358821 $T=54300 36130 0 0 $X=53940 $Y=36000
X776 1 M9_M8_CDNS_7651586358821 $T=57590 18970 0 0 $X=57230 $Y=18840
X777 1 M9_M8_CDNS_7651586358821 $T=57590 27180 0 0 $X=57230 $Y=27050
X778 1 M9_M8_CDNS_7651586358821 $T=58810 43370 0 0 $X=58450 $Y=43240
X779 1 M9_M8_CDNS_7651586358821 $T=74710 18350 0 0 $X=74350 $Y=18220
X780 1 M9_M8_CDNS_7651586358821 $T=74710 26280 0 0 $X=74350 $Y=26150
X781 1 M9_M8_CDNS_7651586358821 $T=74710 34150 0 0 $X=74350 $Y=34020
X782 1 M9_M8_CDNS_7651586358821 $T=74880 9920 0 0 $X=74520 $Y=9790
X783 2 M9_M8_CDNS_7651586358821 $T=77130 16720 0 0 $X=76770 $Y=16590
X784 2 M9_M8_CDNS_7651586358821 $T=77130 24150 0 0 $X=76770 $Y=24020
X785 2 M9_M8_CDNS_7651586358821 $T=77130 33380 0 0 $X=76770 $Y=33250
X786 2 M9_M8_CDNS_7651586358821 $T=78960 40520 0 0 $X=78600 $Y=40390
X787 1 M9_M8_CDNS_7651586358821 $T=83500 11170 0 0 $X=83140 $Y=11040
X788 1 M9_M8_CDNS_7651586358821 $T=85120 19020 0 0 $X=84760 $Y=18890
X789 1 M9_M8_CDNS_7651586358821 $T=85120 28370 0 0 $X=84760 $Y=28240
X790 1 M9_M8_CDNS_7651586358821 $T=85120 35150 0 0 $X=84760 $Y=35020
X791 2 M9_M8_CDNS_7651586358821 $T=99950 62120 0 0 $X=99590 $Y=61990
X792 2 M9_M8_CDNS_7651586358821 $T=100620 51980 0 0 $X=100260 $Y=51850
X793 2 M9_M8_CDNS_7651586358821 $T=102130 14020 0 0 $X=101770 $Y=13890
X794 2 M9_M8_CDNS_7651586358821 $T=102130 22060 0 0 $X=101770 $Y=21930
X795 2 M9_M8_CDNS_7651586358821 $T=102130 29250 0 0 $X=101770 $Y=29120
X796 2 M9_M8_CDNS_7651586358821 $T=102130 38320 0 0 $X=101770 $Y=38190
X797 2 M9_M8_CDNS_7651586358821 $T=105780 67340 0 0 $X=105420 $Y=67210
X798 1 M9_M8_CDNS_7651586358821 $T=106700 9920 0 0 $X=106340 $Y=9790
X799 1 M9_M8_CDNS_7651586358821 $T=106700 18310 0 0 $X=106340 $Y=18180
X800 1 M9_M8_CDNS_7651586358821 $T=106700 26700 0 0 $X=106340 $Y=26570
X801 1 M9_M8_CDNS_7651586358821 $T=106700 35090 0 0 $X=106340 $Y=34960
X802 1 M9_M8_CDNS_7651586358821 $T=106700 46070 0 0 $X=106340 $Y=45940
X803 1 M9_M8_CDNS_7651586358821 $T=106700 55950 0 0 $X=106340 $Y=55820
X804 1 M9_M8_CDNS_7651586358821 $T=106700 61400 0 0 $X=106340 $Y=61270
X805 46 2 1 34 48 47 64 65 142 143 c2mos $T=83140 12860 0 0 $X=83140 $Y=12710
X806 46 2 1 33 49 47 66 67 144 145 c2mos $T=83140 20330 0 0 $X=83140 $Y=20180
X807 46 2 1 35 50 47 68 69 146 147 c2mos $T=83140 29510 0 0 $X=83140 $Y=29360
X808 46 2 1 40 51 47 70 71 148 149 c2mos $T=83140 36740 0 0 $X=83140 $Y=36590
X809 46 2 1 41 52 47 72 73 150 151 c2mos $T=92740 8970 0 0 $X=92740 $Y=8820
X810 46 2 1 9 53 47 74 75 152 153 c2mos $T=92740 16440 0 0 $X=92740 $Y=16290
X811 46 2 1 10 54 47 76 77 154 155 c2mos $T=92740 25620 0 0 $X=92740 $Y=25470
X812 46 2 1 11 55 47 78 79 156 157 c2mos $T=92740 32850 0 0 $X=92740 $Y=32700
X813 46 2 1 8 57 47 80 81 158 159 c2mos $T=98960 56760 0 0 $X=98960 $Y=56610
X814 46 2 1 12 56 47 82 83 160 161 c2mos $T=98990 46730 0 0 $X=98990 $Y=46580
X815 46 2 1 39 58 47 84 85 162 163 c2mos $T=104400 62160 0 0 $X=104400 $Y=62010
X816 3 2 42 1 24 164 86 and2 $T=15650 55370 0 0 $X=12980 $Y=52790
X817 4 2 42 1 39 165 87 and2 $T=15650 65170 0 0 $X=12980 $Y=62590
X818 13 2 42 1 19 166 88 and2 $T=15950 34640 0 0 $X=13280 $Y=32060
X819 14 2 42 1 20 167 89 and2 $T=15950 44110 0 0 $X=13280 $Y=41530
X820 13 2 43 1 15 168 90 and2 $T=24170 29010 0 0 $X=21500 $Y=26430
X821 14 2 43 1 18 169 91 and2 $T=24270 39260 0 0 $X=21600 $Y=36680
X822 3 2 43 1 21 170 92 and2 $T=24270 48510 0 0 $X=21600 $Y=45930
X823 4 2 43 1 23 171 93 and2 $T=24270 58330 0 0 $X=21600 $Y=55750
X824 13 2 44 1 26 172 94 and2 $T=45790 21400 0 0 $X=43120 $Y=18820
X825 14 2 44 1 25 173 95 and2 $T=46640 30040 0 0 $X=43970 $Y=27460
X826 3 2 44 1 28 174 96 and2 $T=47840 38160 0 0 $X=45170 $Y=35580
X827 4 2 44 1 29 175 97 and2 $T=49730 46350 0 0 $X=47060 $Y=43770
X828 13 2 45 1 34 176 98 and2 $T=72230 11810 0 0 $X=69560 $Y=9230
X829 14 2 45 1 33 177 99 and2 $T=72470 21070 0 0 $X=69800 $Y=18490
X830 3 2 45 1 35 178 100 and2 $T=73020 29170 0 0 $X=70350 $Y=26590
X831 4 2 45 1 40 179 101 and2 $T=74450 37230 0 0 $X=71780 $Y=34650
X832 22 15 1 2 5 27 102 half_adder $T=29710 27070 0 0 $X=32010 $Y=27350
X833 23 24 1 2 8 17 104 half_adder $T=30010 51510 0 0 $X=32310 $Y=51790
X834 29 7 1 2 12 31 106 half_adder $T=55120 42950 0 0 $X=57420 $Y=43230
X835 51 55 1 2 59 36 108 half_adder $T=104810 34950 0 0 $X=107110 $Y=35230
X836 18 19 16 2 1 6 22 112 111 113
+ 110 full_adder $T=28640 34740 0 0 $X=30420 $Y=35990
X837 21 20 17 2 1 7 16 116 115 117
+ 114 full_adder $T=28640 43080 0 0 $X=30420 $Y=44330
X838 25 5 30 2 1 10 32 120 119 121
+ 118 full_adder $T=53750 26520 0 0 $X=55530 $Y=27770
X839 28 6 31 2 1 11 30 124 123 125
+ 122 full_adder $T=53750 34740 0 0 $X=55530 $Y=35990
X840 26 27 32 2 1 9 41 128 127 129
+ 126 full_adder $T=54350 18300 0 0 $X=56130 $Y=19550
X841 50 54 36 2 1 60 38 132 131 133
+ 130 full_adder $T=104430 26180 0 0 $X=106210 $Y=27430
X842 49 53 38 2 1 61 37 136 135 137
+ 134 full_adder $T=105090 17720 0 0 $X=106870 $Y=18970
X843 48 52 37 2 1 62 63 140 139 141
+ 138 full_adder $T=105100 9270 0 0 $X=106880 $Y=10520
M0 64 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=83890 $Y=13510 $dt=0
M1 66 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=83890 $Y=20980 $dt=0
M2 68 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=83890 $Y=30160 $dt=0
M3 70 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=83890 $Y=37390 $dt=0
M4 1 47 48 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=91350 $Y=13030 $dt=0
M5 1 47 49 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=91350 $Y=20500 $dt=0
M6 1 47 50 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=91350 $Y=29680 $dt=0
M7 1 47 51 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=91350 $Y=36910 $dt=0
M8 72 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=93490 $Y=9620 $dt=0
M9 74 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=93490 $Y=17090 $dt=0
M10 76 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=93490 $Y=26270 $dt=0
M11 78 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=93490 $Y=33500 $dt=0
M12 80 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=99710 $Y=57410 $dt=0
M13 82 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=99740 $Y=47380 $dt=0
M14 1 47 52 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=100950 $Y=9140 $dt=0
M15 1 47 53 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=100950 $Y=16610 $dt=0
M16 1 47 54 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=100950 $Y=25790 $dt=0
M17 1 47 55 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=100950 $Y=33020 $dt=0
M18 84 46 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.48209 scb=0.00151892 scc=4.69814e-06 $X=105150 $Y=62810 $dt=0
M19 1 47 57 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=107170 $Y=56930 $dt=0
M20 1 47 56 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=107200 $Y=46900 $dt=0
M21 1 47 58 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=112610 $Y=62330 $dt=0
M22 86 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=13400 $Y=56300 $dt=1
M23 87 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=13400 $Y=66100 $dt=1
M24 88 13 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=13700 $Y=35570 $dt=1
M25 89 14 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=13700 $Y=45040 $dt=1
M26 2 3 86 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=13810 $Y=56300 $dt=1
M27 2 4 87 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=13810 $Y=66100 $dt=1
M28 2 13 88 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=14110 $Y=35570 $dt=1
M29 2 14 89 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=14110 $Y=45040 $dt=1
M30 86 42 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=14700 $Y=56300 $dt=1
M31 87 42 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=14700 $Y=66100 $dt=1
M32 88 42 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=15000 $Y=35570 $dt=1
M33 89 42 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=15000 $Y=45040 $dt=1
M34 90 13 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=21920 $Y=29940 $dt=1
M35 91 14 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=22020 $Y=40190 $dt=1
M36 92 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=22020 $Y=49440 $dt=1
M37 93 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=22020 $Y=59260 $dt=1
M38 2 13 90 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=22330 $Y=29940 $dt=1
M39 2 14 91 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=22430 $Y=40190 $dt=1
M40 2 3 92 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=22430 $Y=49440 $dt=1
M41 2 4 93 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=22430 $Y=59260 $dt=1
M42 90 43 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=23220 $Y=29940 $dt=1
M43 91 43 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=23320 $Y=40190 $dt=1
M44 92 43 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=23320 $Y=49440 $dt=1
M45 93 43 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=23320 $Y=59260 $dt=1
M46 94 13 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=43540 $Y=22330 $dt=1
M47 2 13 94 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=43950 $Y=22330 $dt=1
M48 95 14 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=44390 $Y=30970 $dt=1
M49 2 14 95 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=44800 $Y=30970 $dt=1
M50 94 44 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=44840 $Y=22330 $dt=1
M51 96 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=45590 $Y=39090 $dt=1
M52 95 44 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=45690 $Y=30970 $dt=1
M53 2 3 96 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=46000 $Y=39090 $dt=1
M54 96 44 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=46890 $Y=39090 $dt=1
M55 97 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=47480 $Y=47280 $dt=1
M56 2 4 97 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=47890 $Y=47280 $dt=1
M57 97 44 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=48780 $Y=47280 $dt=1
M58 98 13 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=69980 $Y=12740 $dt=1
M59 99 14 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=70220 $Y=22000 $dt=1
M60 2 13 98 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=70390 $Y=12740 $dt=1
M61 2 14 99 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=70630 $Y=22000 $dt=1
M62 100 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=70770 $Y=30100 $dt=1
M63 2 3 100 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=71180 $Y=30100 $dt=1
M64 98 45 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=71280 $Y=12740 $dt=1
M65 99 45 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=71520 $Y=22000 $dt=1
M66 100 45 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=72070 $Y=30100 $dt=1
M67 101 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=72200 $Y=38160 $dt=1
M68 2 4 101 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=72610 $Y=38160 $dt=1
M69 101 45 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=73500 $Y=38160 $dt=1
.ends pipeline_mult
