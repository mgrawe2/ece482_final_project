* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mult_auto                                    *
* Netlisted  : Sat Dec  6 18:47:50 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765068464210                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765068464210 S_source_0 S_source_2 D_drain_1 4 5
** N=5 EP=5 FDC=2
M0 D_drain_1 4 S_source_0 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 S_source_2 4 D_drain_1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765068464210

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765068464212                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765068464212 S_source_0 D_drain_1 3 S_source_2 5
** N=5 EP=5 FDC=2
M0 D_drain_1 3 S_source_0 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 S_source_2 3 D_drain_1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765068464212

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv IN VDD OUT VSS
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X4 VSS OUT IN VSS VSS nmos1v_CDNS_765068464212 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 A VDD B VSS OUT 7
*.DEVICECLIMB
** N=7 EP=6 FDC=9
X10 6 6 7 A VSS nmos1v_CDNS_765068464210 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 6 6 VSS B VSS nmos1v_CDNS_765068464210 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X14 7 VDD OUT VSS inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 VDD B 7 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M1 OUT 7 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M2 VDD 7 OUT VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor B VDD VSS B_bar OUT A
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X8 OUT A B_bar OUT VSS nmos1v_CDNS_765068464212 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X9 B_bar OUT A B_bar VSS nmos1v_CDNS_765068464212 $T=800 -1920 0 0 $X=380 $Y=-2120
X10 B VDD B_bar VSS inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
M0 OUT B A VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 OUT A B VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 B A OUT VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder B A VSS VDD S Co
** N=9 EP=6 FDC=24
X6 A VDD B VSS Co 8 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X10 B VDD VSS 7 S A xor $T=4660 3560 0 0 $X=2440 $Y=1000
M0 7 B VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2860 $Y=3790 $dt=1
M1 VDD B 7 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3270 $Y=3790 $dt=1
M2 A B S VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4160 $Y=3790 $dt=1
M3 8 A VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6760 $Y=3790 $dt=1
M4 VDD A 8 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7170 $Y=3790 $dt=1
M5 8 B VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8060 $Y=3790 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765068464213                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765068464213 S_source_0 D_drain_1 3 S_source_2 D_drain_3 6 7 S_source_4 9
** N=9 EP=9 FDC=4
M0 D_drain_1 3 S_source_0 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 S_source_2 6 D_drain_1 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 D_drain_3 7 S_source_2 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 S_source_4 9 D_drain_3 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_765068464213

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765068464214                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765068464214 S_source_0 D_drain_1 S_source_2 4 5 D_drain_3 S_source_4 8 9 B
** N=11 EP=10 FDC=4
M0 D_drain_1 4 S_source_0 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 S_source_2 5 D_drain_1 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 D_drain_3 8 S_source_2 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 S_source_4 9 D_drain_3 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_765068464214

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network OUT P Ci VDD VSS P_bar A
** N=11 EP=7 FDC=8
X12 OUT 8 Ci VSS 9 P P_bar OUT A nmos1v_CDNS_765068464213 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 OUT 10 VDD Ci P_bar 11 OUT P A VDD pmos1v_CDNS_765068464214 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder B A Ci VDD VSS S Co
** N=15 EP=7 FDC=36
X14 10 VDD Co VSS inv $T=12350 3410 0 0 $X=11870 $Y=1250
X19 B VDD VSS 11 9 A xor $T=4170 3810 0 0 $X=1950 $Y=1250
X20 9 VDD VSS 8 S Ci xor $T=8070 3810 0 0 $X=5850 $Y=1250
X23 10 9 Ci VDD VSS 8 A fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 11 B VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 VDD B 11 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 A B 9 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 8 9 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 VDD 9 8 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 Ci 9 S VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 Co 10 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 VDD 10 Co VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mult_auto                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mult_auto A0 A1 A2 A3 B0 B1 B2 B3 P0 P1
+ P2 P3 P4 P5 P6 P7 VDD VSS
** N=143 EP=18 FDC=576
X584 A1 VDD B0 VSS 3 52 and2 $T=5890 68510 0 0 $X=3220 $Y=65930
X585 A0 VDD B0 VSS P0 53 and2 $T=5890 78310 0 0 $X=3220 $Y=75730
X586 A3 VDD B0 VSS 5 54 and2 $T=6190 47780 0 0 $X=3520 $Y=45200
X587 A2 VDD B0 VSS 6 55 and2 $T=6190 57250 0 0 $X=3520 $Y=54670
X588 A3 VDD B1 VSS 7 56 and2 $T=14410 42150 0 0 $X=11740 $Y=39570
X589 A2 VDD B1 VSS 10 57 and2 $T=14510 52400 0 0 $X=11840 $Y=49820
X590 A1 VDD B1 VSS 8 58 and2 $T=14510 61650 0 0 $X=11840 $Y=59070
X591 A0 VDD B1 VSS 9 59 and2 $T=14510 71470 0 0 $X=11840 $Y=68890
X592 A3 VDD B2 VSS 11 60 and2 $T=36030 34540 0 0 $X=33360 $Y=31960
X593 A2 VDD B2 VSS 12 61 and2 $T=36880 43180 0 0 $X=34210 $Y=40600
X594 A1 VDD B2 VSS 13 62 and2 $T=38080 51300 0 0 $X=35410 $Y=48720
X595 A0 VDD B2 VSS 14 63 and2 $T=39970 59490 0 0 $X=37300 $Y=56910
X596 A3 VDD B3 VSS 15 64 and2 $T=62470 24950 0 0 $X=59800 $Y=22370
X597 A2 VDD B3 VSS 16 65 and2 $T=62710 34210 0 0 $X=60040 $Y=31630
X598 A1 VDD B3 VSS 17 66 and2 $T=63260 42310 0 0 $X=60590 $Y=39730
X599 A0 VDD B3 VSS 18 67 and2 $T=64690 50370 0 0 $X=62020 $Y=47790
X600 38 7 VSS VDD 29 39 half_adder $T=19950 40210 0 0 $X=22250 $Y=40490
X601 9 3 VSS VDD P1 37 half_adder $T=20250 64650 0 0 $X=22550 $Y=64930
X602 14 31 VSS VDD P2 41 half_adder $T=45360 56090 0 0 $X=47660 $Y=56370
X603 18 34 VSS VDD P3 44 half_adder $T=69570 48090 0 0 $X=71870 $Y=48370
X604 10 5 36 VDD VSS 30 38 full_adder $T=18880 47880 0 0 $X=20660 $Y=49130
X605 8 6 37 VDD VSS 31 36 full_adder $T=18880 56220 0 0 $X=20660 $Y=57470
X606 12 29 40 VDD VSS 33 42 full_adder $T=43990 39660 0 0 $X=45770 $Y=40910
X607 13 30 41 VDD VSS 34 40 full_adder $T=43990 47880 0 0 $X=45770 $Y=49130
X608 11 39 42 VDD VSS 32 43 full_adder $T=44590 31440 0 0 $X=46370 $Y=32690
X609 17 33 44 VDD VSS P4 46 full_adder $T=69190 39320 0 0 $X=70970 $Y=40570
X610 16 32 46 VDD VSS P5 45 full_adder $T=69850 30860 0 0 $X=71630 $Y=32110
X611 15 43 45 VDD VSS P6 P7 full_adder $T=69860 22410 0 0 $X=71640 $Y=23660
M0 52 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3640 $Y=69440 $dt=1
M1 53 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3640 $Y=79240 $dt=1
M2 54 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3940 $Y=48710 $dt=1
M3 55 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3940 $Y=58180 $dt=1
M4 VDD A1 52 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4050 $Y=69440 $dt=1
M5 VDD A0 53 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4050 $Y=79240 $dt=1
M6 VDD A3 54 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4350 $Y=48710 $dt=1
M7 VDD A2 55 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4350 $Y=58180 $dt=1
M8 52 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4940 $Y=69440 $dt=1
M9 53 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4940 $Y=79240 $dt=1
M10 54 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=5240 $Y=48710 $dt=1
M11 55 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=5240 $Y=58180 $dt=1
M12 56 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12160 $Y=43080 $dt=1
M13 57 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=53330 $dt=1
M14 58 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=62580 $dt=1
M15 59 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=72400 $dt=1
M16 VDD A3 56 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12570 $Y=43080 $dt=1
M17 VDD A2 57 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=53330 $dt=1
M18 VDD A1 58 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=62580 $dt=1
M19 VDD A0 59 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=72400 $dt=1
M20 56 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13460 $Y=43080 $dt=1
M21 57 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=53330 $dt=1
M22 58 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=62580 $dt=1
M23 59 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=72400 $dt=1
M24 60 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=33780 $Y=35470 $dt=1
M25 VDD A3 60 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=34190 $Y=35470 $dt=1
M26 61 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=34630 $Y=44110 $dt=1
M27 VDD A2 61 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=35040 $Y=44110 $dt=1
M28 60 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=35080 $Y=35470 $dt=1
M29 62 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=35830 $Y=52230 $dt=1
M30 61 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=35930 $Y=44110 $dt=1
M31 VDD A1 62 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=36240 $Y=52230 $dt=1
M32 62 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=37130 $Y=52230 $dt=1
M33 63 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=37720 $Y=60420 $dt=1
M34 VDD A0 63 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=38130 $Y=60420 $dt=1
M35 63 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=39020 $Y=60420 $dt=1
M36 64 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=60220 $Y=25880 $dt=1
M37 65 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=60460 $Y=35140 $dt=1
M38 VDD A3 64 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=60630 $Y=25880 $dt=1
M39 VDD A2 65 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=60870 $Y=35140 $dt=1
M40 66 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=61010 $Y=43240 $dt=1
M41 VDD A1 66 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=61420 $Y=43240 $dt=1
M42 64 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=61520 $Y=25880 $dt=1
M43 65 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=61760 $Y=35140 $dt=1
M44 66 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=62310 $Y=43240 $dt=1
M45 67 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=62440 $Y=51300 $dt=1
M46 VDD A0 67 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=62850 $Y=51300 $dt=1
M47 67 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=63740 $Y=51300 $dt=1
.ends mult_auto
