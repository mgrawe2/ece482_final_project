* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : fa_co_network                                *
* Netlisted  : Thu Dec  4 13:03:23 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764874998100                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764874998100 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764874998100

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764874998101                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764874998101 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764874998101

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764874998104                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764874998104 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764874998104

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764874998100                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764874998100 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_764874998100

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764874998101                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764874998101 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=45.4346 scb=0.0376748 scc=0.00495816 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=31.5894 scb=0.0205288 scc=0.00239824 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=31.5894 scb=0.0205288 scc=0.00239824 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=45.4346 scb=0.0376748 scc=0.00495816 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_764874998101

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 5 4 3 1 2 10 7
** N=11 EP=7 FDC=8
X0 1 M1_PO_CDNS_764874998100 $T=-220 -60 0 0 $X=-320 $Y=-180
X1 2 M1_PO_CDNS_764874998100 $T=-210 730 0 0 $X=-310 $Y=610
X2 2 M1_PO_CDNS_764874998100 $T=190 -60 0 0 $X=90 $Y=-180
X3 1 M1_PO_CDNS_764874998100 $T=200 730 0 0 $X=100 $Y=610
X4 3 M2_M1_CDNS_764874998101 $T=-830 -970 0 0 $X=-910 $Y=-1100
X5 1 M2_M1_CDNS_764874998101 $T=-220 -60 0 0 $X=-300 $Y=-190
X6 1 M2_M1_CDNS_764874998101 $T=200 730 0 0 $X=120 $Y=600
X7 3 M2_M1_CDNS_764874998101 $T=810 -970 0 0 $X=730 $Y=-1100
X8 4 M1_PO_CDNS_764874998104 $T=-590 550 0 0 $X=-690 $Y=190
X9 5 M1_PO_CDNS_764874998104 $T=570 550 0 0 $X=470 $Y=190
X10 3 6 4 7 8 1 2 3 5 nmos1v_CDNS_764874998100 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X11 3 9 10 4 2 11 3 1 5 7
+ 10 pmos1v_CDNS_764874998101 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network
