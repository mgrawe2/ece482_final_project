* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : full_adder                                   *
* Netlisted  : Thu Dec  4 16:56:35 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_764888989950                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_764888989950 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_764888989950

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764888989951                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764888989951 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764888989951

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764888989952                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764888989952 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764888989952

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888989953                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888989953 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888989953

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888989954                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888989954 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888989954

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888989955                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888989955 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888989955

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_7648889899512                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_7648889899512 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_7648889899512

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7648889899513                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7648889899513 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7648889899513

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_7648889899514                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_7648889899514 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_7648889899514

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764888989950                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764888989950 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_764888989950

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764888989951                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764888989951 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764888989951

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X0 2 M1_NWELL_CDNS_7648889899512 $T=190 2570 0 0 $X=-230 $Y=2270
X1 1 M1_PO_CDNS_7648889899513 $T=-160 30 0 0 $X=-260 $Y=-330
X2 4 M1_PSUB_CDNS_7648889899514 $T=190 -2020 0 0 $X=-190 $Y=-2160
X3 2 3 1 2 4 2 pmos1v_CDNS_764888989950 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 3 1 4 4 nmos1v_CDNS_764888989951 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888989957                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888989957 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888989957

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764888989959                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764888989959 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764888989959

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X0 6 M2_M1_CDNS_764888989953 $T=-30 -450 0 0 $X=-160 $Y=-580
X1 5 M2_M1_CDNS_764888989953 $T=1330 -190 0 0 $X=1200 $Y=-320
X2 6 M2_M1_CDNS_764888989954 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X3 6 M2_M1_CDNS_764888989954 $T=-250 380 0 0 $X=-380 $Y=250
X4 5 M2_M1_CDNS_764888989957 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X5 5 M2_M1_CDNS_764888989957 $T=-660 950 0 0 $X=-740 $Y=700
X6 5 M2_M1_CDNS_764888989957 $T=160 -1560 0 0 $X=80 $Y=-1810
X7 5 M2_M1_CDNS_764888989957 $T=160 950 0 0 $X=80 $Y=700
X8 5 M2_M1_CDNS_764888989957 $T=1050 -1560 0 0 $X=970 $Y=-1810
X9 5 M2_M1_CDNS_764888989957 $T=1050 950 0 0 $X=970 $Y=700
X10 1 M1_PO_CDNS_764888989959 $T=-450 10 0 0 $X=-550 $Y=-110
X11 1 M1_PO_CDNS_764888989959 $T=-450 1890 0 0 $X=-550 $Y=1770
X12 3 M1_PO_CDNS_764888989959 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X13 1 M1_PO_CDNS_764888989959 $T=-40 1890 0 0 $X=-140 $Y=1770
X14 6 M1_PO_CDNS_764888989959 $T=850 -980 0 0 $X=750 $Y=-1100
X15 5 6 1 5 4 2 pmos1v_CDNS_764888989950 $T=-500 230 0 0 $X=-920 $Y=30
X16 1 5 6 1 4 2 pmos1v_CDNS_764888989950 $T=800 230 0 0 $X=380 $Y=30
X17 5 6 3 5 4 nmos1v_CDNS_764888989951 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X18 3 5 6 3 4 nmos1v_CDNS_764888989951 $T=800 -1920 0 0 $X=380 $Y=-2120
X19 1 2 3 4 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
M0 5 1 6 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 5 6 1 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 1 6 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764888989952                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764888989952 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_764888989952

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764888989953                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764888989953 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_764888989953

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=8
X0 1 M2_M1_CDNS_764888989955 $T=-830 -970 0 0 $X=-910 $Y=-1100
X1 2 M2_M1_CDNS_764888989955 $T=-220 -60 0 0 $X=-300 $Y=-190
X2 2 M2_M1_CDNS_764888989955 $T=200 730 0 0 $X=120 $Y=600
X3 1 M2_M1_CDNS_764888989955 $T=810 -970 0 0 $X=730 $Y=-1100
X4 2 M1_PO_CDNS_764888989959 $T=-220 -60 0 0 $X=-320 $Y=-180
X5 5 M1_PO_CDNS_764888989959 $T=-210 730 0 0 $X=-310 $Y=610
X6 5 M1_PO_CDNS_764888989959 $T=190 -60 0 0 $X=90 $Y=-180
X7 2 M1_PO_CDNS_764888989959 $T=200 730 0 0 $X=100 $Y=610
X8 4 M1_NWELL_CDNS_7648889899512 $T=-10 2990 0 0 $X=-430 $Y=2690
X9 3 M1_PO_CDNS_7648889899513 $T=-590 550 0 0 $X=-690 $Y=190
X10 7 M1_PO_CDNS_7648889899513 $T=570 550 0 0 $X=470 $Y=190
X11 6 M1_PSUB_CDNS_7648889899514 $T=0 -1600 0 0 $X=-380 $Y=-1740
X12 1 8 3 6 9 2 5 1 7 nmos1v_CDNS_764888989952 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 1 10 4 3 5 11 1 2 7 6
+ 4 pmos1v_CDNS_764888989953 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 1 2 5 4 3 6 10
** N=15 EP=7 FDC=36
X0 1 M4_M3_CDNS_764888989950 $T=6980 3080 0 0 $X=6900 $Y=2950
X1 1 M4_M3_CDNS_764888989950 $T=10140 2970 0 0 $X=10060 $Y=2840
X2 2 M3_M2_CDNS_764888989951 $T=2270 3860 0 0 $X=2190 $Y=3730
X3 1 M3_M2_CDNS_764888989951 $T=5790 3080 0 0 $X=5710 $Y=2950
X4 3 M3_M2_CDNS_764888989951 $T=9120 4760 0 0 $X=9040 $Y=4630
X5 1 M3_M2_CDNS_764888989951 $T=11410 2940 0 0 $X=11330 $Y=2810
X6 4 M3_M2_CDNS_764888989951 $T=12920 3510 0 0 $X=12840 $Y=3380
X7 5 M3_M2_CDNS_764888989952 $T=7300 3360 0 0 $X=7170 $Y=3230
X8 5 M3_M2_CDNS_764888989952 $T=10110 3640 0 0 $X=9980 $Y=3510
X9 6 M2_M1_CDNS_764888989953 $T=6470 5920 0 0 $X=6340 $Y=5790
X10 5 M2_M1_CDNS_764888989953 $T=7620 3360 0 0 $X=7490 $Y=3230
X11 5 M2_M1_CDNS_764888989953 $T=10320 3640 0 0 $X=10190 $Y=3510
X12 6 M2_M1_CDNS_764888989954 $T=3420 5920 0 0 $X=3290 $Y=5790
X13 1 M2_M1_CDNS_764888989955 $T=5250 3070 0 0 $X=5170 $Y=2940
X14 7 M2_M1_CDNS_764888989955 $T=9530 2380 0 0 $X=9450 $Y=2250
X15 8 M2_M1_CDNS_764888989955 $T=9530 5090 0 0 $X=9450 $Y=4960
X16 6 M2_M1_CDNS_764888989955 $T=10820 5970 0 0 $X=10740 $Y=5840
X17 7 M2_M1_CDNS_764888989955 $T=11040 2940 0 0 $X=10960 $Y=2810
X18 1 M2_M1_CDNS_764888989955 $T=11390 3320 0 0 $X=11310 $Y=3190
X19 4 M2_M1_CDNS_764888989955 $T=12920 3510 0 0 $X=12840 $Y=3380
X20 9 6 4 10 inv $T=12350 3410 0 0 $X=11870 $Y=1250
X21 2 6 11 10 8 1 xor $T=4170 3810 0 0 $X=1950 $Y=1250
X22 8 6 7 10 3 5 xor $T=8070 3810 0 0 $X=5850 $Y=1250
X23 9 8 5 6 7 10 1 12 13 14
+ 15 fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 11 2 6 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 6 2 11 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 1 2 8 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 7 8 6 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 6 8 7 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 5 8 3 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 4 9 6 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 6 9 4 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder
