* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : and2_auto                                    *
* Netlisted  : Wed Dec  3 21:39:32 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764819567080                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764819567080 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_764819567080

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764819567081                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764819567081 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764819567081

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_764819567082                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_764819567082 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_764819567082

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764819567083                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764819567083 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764819567083

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764819567080                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764819567080 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764819567080

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764819567081                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764819567081 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_764819567081

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764819567082                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764819567082 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 4 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 3 4 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764819567082

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
** N=4 EP=4 FDC=4
X0 1 M1_NWELL_CDNS_764819567080 $T=190 2570 0 0 $X=-230 $Y=2270
X1 2 M1_PSUB_CDNS_764819567082 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 3 M1_PO_CDNS_764819567083 $T=-160 30 0 0 $X=-260 $Y=-330
X3 4 1 1 3 2 1 pmos1v_CDNS_764819567081 $T=-60 630 0 0 $X=-480 $Y=430
X4 2 4 2 3 2 nmos1v_CDNS_764819567082 $T=-60 -1520 0 0 $X=-480 $Y=-1720
M0 4 3 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-60 $Y=630 $dt=1
M1 1 3 4 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=350 $Y=630 $dt=1
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2_auto                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2_auto 5 6 7 1 4
** N=7 EP=5 FDC=12
X0 1 M1_NWELL_CDNS_764819567080 $T=3500 8780 0 0 $X=3080 $Y=8480
X1 2 M2_M1_CDNS_764819567081 $T=2440 4690 0 0 $X=2360 $Y=4440
X2 3 M2_M1_CDNS_764819567081 $T=2850 7560 0 0 $X=2770 $Y=7310
X3 2 M2_M1_CDNS_764819567081 $T=3260 4690 0 0 $X=3180 $Y=4440
X4 2 M2_M1_CDNS_764819567081 $T=3740 4690 0 0 $X=3660 $Y=4440
X5 3 M2_M1_CDNS_764819567081 $T=4150 7560 0 0 $X=4070 $Y=7310
X6 2 M2_M1_CDNS_764819567081 $T=4560 4690 0 0 $X=4480 $Y=4440
X7 4 M1_PSUB_CDNS_764819567082 $T=4150 3470 0 0 $X=3770 $Y=3330
X8 5 M1_PO_CDNS_764819567083 $T=2500 6270 0 0 $X=2400 $Y=5910
X9 6 M1_PO_CDNS_764819567083 $T=3800 5970 0 0 $X=3700 $Y=5610
X10 2 2 3 5 4 nmos1v_CDNS_764819567080 $T=2600 3970 0 0 $X=2180 $Y=3770
X11 2 2 4 6 4 nmos1v_CDNS_764819567080 $T=3900 3970 0 0 $X=3480 $Y=3770
X12 3 1 1 5 4 1 pmos1v_CDNS_764819567081 $T=2600 6840 0 0 $X=2180 $Y=6640
X13 3 1 1 6 4 1 pmos1v_CDNS_764819567081 $T=3900 6840 0 0 $X=3480 $Y=6640
X14 1 4 3 7 inv $T=5260 6210 0 0 $X=4780 $Y=4050
M0 3 5 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2600 $Y=6840 $dt=1
M1 1 5 3 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3010 $Y=6840 $dt=1
M2 3 6 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3900 $Y=6840 $dt=1
M3 1 6 3 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4310 $Y=6840 $dt=1
.ends and2_auto
