* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mult_auto                                    *
* Netlisted  : Sat Dec  6 15:35:26 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765056920380                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765056920380 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765056920380

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765056920381                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765056920381 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765056920381

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765056920382                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765056920382 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765056920382

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765056920383                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765056920383 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765056920383

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765056920384                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765056920384 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765056920384

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765056920385                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765056920385 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765056920385

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765056920386                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765056920386 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765056920386

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765056920387                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765056920387 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765056920387

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765056920388                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765056920388 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765056920388

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_7650569203810                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_7650569203810 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_7650569203810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7650569203811                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7650569203811 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7650569203811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_7650569203812                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_7650569203812 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_7650569203812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7650569203813                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7650569203813 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7650569203813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765056920380                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765056920380 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765056920380

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765056920381                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765056920381 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_765056920381

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765056920382                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765056920382 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765056920382

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=2
X0 2 M1_NWELL_CDNS_7650569203810 $T=190 2570 0 0 $X=-230 $Y=2270
X1 4 M1_PSUB_CDNS_7650569203812 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 1 M1_PO_CDNS_7650569203813 $T=-160 30 0 0 $X=-260 $Y=-330
X3 2 3 1 2 5 2 pmos1v_CDNS_765056920381 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 3 1 4 5 nmos1v_CDNS_765056920382 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7 8
*.DEVICECLIMB
** N=8 EP=8 FDC=9
X0 2 M1_NWELL_CDNS_7650569203810 $T=-1350 2870 0 0 $X=-1770 $Y=2570
X1 7 M2_M1_CDNS_7650569203811 $T=-2410 -1220 0 0 $X=-2490 $Y=-1470
X2 8 M2_M1_CDNS_7650569203811 $T=-2000 1650 0 0 $X=-2080 $Y=1400
X3 7 M2_M1_CDNS_7650569203811 $T=-1590 -1220 0 0 $X=-1670 $Y=-1470
X4 7 M2_M1_CDNS_7650569203811 $T=-1110 -1220 0 0 $X=-1190 $Y=-1470
X5 8 M2_M1_CDNS_7650569203811 $T=-700 1650 0 0 $X=-780 $Y=1400
X6 7 M2_M1_CDNS_7650569203811 $T=-290 -1220 0 0 $X=-370 $Y=-1470
X7 4 M1_PSUB_CDNS_7650569203812 $T=-700 -2440 0 0 $X=-1080 $Y=-2580
X8 1 M1_PO_CDNS_7650569203813 $T=-2350 360 0 0 $X=-2450 $Y=0
X9 3 M1_PO_CDNS_7650569203813 $T=-1050 60 0 0 $X=-1150 $Y=-300
X10 7 7 8 1 6 nmos1v_CDNS_765056920380 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 7 7 4 3 6 nmos1v_CDNS_765056920380 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X12 2 8 1 2 6 2 pmos1v_CDNS_765056920381 $T=-2250 930 0 0 $X=-2670 $Y=730
X13 2 8 3 2 6 2 pmos1v_CDNS_765056920381 $T=-950 930 0 0 $X=-1370 $Y=730
X14 8 2 5 4 6 inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 2 3 8 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M1 5 8 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M2 2 8 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7650569203814                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7650569203814 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7650569203814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7650569203815                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7650569203815 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7650569203815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7650569203818                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7650569203818 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7650569203818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=9
X0 5 M2_M1_CDNS_7650569203811 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X1 5 M2_M1_CDNS_7650569203811 $T=-660 950 0 0 $X=-740 $Y=700
X2 5 M2_M1_CDNS_7650569203811 $T=160 -1560 0 0 $X=80 $Y=-1810
X3 5 M2_M1_CDNS_7650569203811 $T=160 950 0 0 $X=80 $Y=700
X4 5 M2_M1_CDNS_7650569203811 $T=1050 -1560 0 0 $X=970 $Y=-1810
X5 5 M2_M1_CDNS_7650569203811 $T=1050 950 0 0 $X=970 $Y=700
X6 5 6 1 5 7 2 pmos1v_CDNS_765056920381 $T=-500 230 0 0 $X=-920 $Y=30
X7 1 5 6 1 7 2 pmos1v_CDNS_765056920381 $T=800 230 0 0 $X=380 $Y=30
X8 5 6 3 5 7 nmos1v_CDNS_765056920382 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X9 3 5 6 3 7 nmos1v_CDNS_765056920382 $T=800 -1920 0 0 $X=380 $Y=-2120
X10 1 2 3 4 7 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
X11 6 M2_M1_CDNS_7650569203814 $T=-30 -450 0 0 $X=-160 $Y=-580
X12 5 M2_M1_CDNS_7650569203814 $T=1330 -190 0 0 $X=1200 $Y=-320
X13 6 M2_M1_CDNS_7650569203815 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X14 6 M2_M1_CDNS_7650569203815 $T=-250 380 0 0 $X=-380 $Y=250
X15 1 M1_PO_CDNS_7650569203818 $T=-450 10 0 0 $X=-550 $Y=-110
X16 1 M1_PO_CDNS_7650569203818 $T=-450 1890 0 0 $X=-550 $Y=1770
X17 3 M1_PO_CDNS_7650569203818 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X18 1 M1_PO_CDNS_7650569203818 $T=-40 1890 0 0 $X=-140 $Y=1770
X19 6 M1_PO_CDNS_7650569203818 $T=850 -980 0 0 $X=750 $Y=-1100
M0 5 1 6 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 5 6 1 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 1 6 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 7 8
** N=10 EP=8 FDC=24
X0 6 M2_M1_CDNS_765056920381 $T=9970 3310 0 0 $X=9890 $Y=3180
X1 5 M2_M1_CDNS_765056920381 $T=10180 2730 0 0 $X=10100 $Y=2600
X2 1 M3_M2_CDNS_765056920388 $T=2760 3570 0 0 $X=2680 $Y=3440
X3 2 M3_M2_CDNS_765056920388 $T=4630 3110 0 0 $X=4550 $Y=2980
X4 6 M3_M2_CDNS_765056920388 $T=9970 3310 0 0 $X=9890 $Y=3180
X5 5 M3_M2_CDNS_765056920388 $T=10180 2730 0 0 $X=10100 $Y=2600
X6 2 3 1 4 6 7 10 9 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X7 1 M2_M1_CDNS_7650569203814 $T=2760 2580 0 0 $X=2630 $Y=2450
X8 1 M2_M1_CDNS_7650569203814 $T=7960 2810 0 0 $X=7830 $Y=2680
X9 5 M2_M1_CDNS_7650569203815 $T=6360 3430 0 0 $X=6230 $Y=3300
X10 1 3 8 4 5 2 7 xor $T=4660 3560 0 0 $X=2440 $Y=1000
M0 8 1 3 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2860 $Y=3790 $dt=1
M1 3 1 8 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3270 $Y=3790 $dt=1
M2 2 1 5 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4160 $Y=3790 $dt=1
M3 9 2 3 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6760 $Y=3790 $dt=1
M4 3 2 9 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7170 $Y=3790 $dt=1
M5 9 1 3 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8060 $Y=3790 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7650569203821                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7650569203821 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7650569203821

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765056920383                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765056920383 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 FDC=4
M0 2 3 1 10 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 10 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 10 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 10 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_765056920383

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765056920384                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765056920384 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_765056920384

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=8
X0 1 M2_M1_CDNS_765056920381 $T=-830 -970 0 0 $X=-910 $Y=-1100
X1 2 M2_M1_CDNS_765056920381 $T=-220 -60 0 0 $X=-300 $Y=-190
X2 2 M2_M1_CDNS_765056920381 $T=200 730 0 0 $X=120 $Y=600
X3 1 M2_M1_CDNS_765056920381 $T=810 -970 0 0 $X=730 $Y=-1100
X4 4 M1_NWELL_CDNS_7650569203810 $T=-10 2990 0 0 $X=-430 $Y=2690
X5 5 M1_PSUB_CDNS_7650569203812 $T=0 -1600 0 0 $X=-380 $Y=-1740
X6 3 M1_PO_CDNS_7650569203813 $T=-590 550 0 0 $X=-690 $Y=190
X7 7 M1_PO_CDNS_7650569203813 $T=570 550 0 0 $X=470 $Y=190
X8 2 M1_PO_CDNS_7650569203818 $T=-220 -60 0 0 $X=-320 $Y=-180
X9 6 M1_PO_CDNS_7650569203818 $T=-210 730 0 0 $X=-310 $Y=610
X10 6 M1_PO_CDNS_7650569203818 $T=190 -60 0 0 $X=90 $Y=-180
X11 2 M1_PO_CDNS_7650569203818 $T=200 730 0 0 $X=100 $Y=610
X12 1 9 3 5 10 2 6 1 7 8 nmos1v_CDNS_765056920383 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 1 11 4 3 6 12 1 2 7 8
+ 4 pmos1v_CDNS_765056920384 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=16 EP=12 FDC=36
X0 2 M2_M1_CDNS_765056920381 $T=5250 3070 0 0 $X=5170 $Y=2940
X1 9 M2_M1_CDNS_765056920381 $T=9530 2380 0 0 $X=9450 $Y=2250
X2 10 M2_M1_CDNS_765056920381 $T=9530 5090 0 0 $X=9450 $Y=4960
X3 4 M2_M1_CDNS_765056920381 $T=10820 5970 0 0 $X=10740 $Y=5840
X4 9 M2_M1_CDNS_765056920381 $T=11040 2940 0 0 $X=10960 $Y=2810
X5 2 M2_M1_CDNS_765056920381 $T=11390 3320 0 0 $X=11310 $Y=3190
X6 7 M2_M1_CDNS_765056920381 $T=12920 3510 0 0 $X=12840 $Y=3380
X7 2 M4_M3_CDNS_765056920387 $T=6980 3080 0 0 $X=6900 $Y=2950
X8 2 M4_M3_CDNS_765056920387 $T=10140 2970 0 0 $X=10060 $Y=2840
X9 1 M3_M2_CDNS_765056920388 $T=2270 3860 0 0 $X=2190 $Y=3730
X10 2 M3_M2_CDNS_765056920388 $T=5790 3080 0 0 $X=5710 $Y=2950
X11 6 M3_M2_CDNS_765056920388 $T=9120 4760 0 0 $X=9040 $Y=4630
X12 2 M3_M2_CDNS_765056920388 $T=11410 2940 0 0 $X=11330 $Y=2810
X13 7 M3_M2_CDNS_765056920388 $T=12920 3510 0 0 $X=12840 $Y=3380
X14 11 4 7 5 8 inv $T=12350 3410 0 0 $X=11870 $Y=1250
X15 4 M2_M1_CDNS_7650569203814 $T=6470 5920 0 0 $X=6340 $Y=5790
X16 3 M2_M1_CDNS_7650569203814 $T=7620 3360 0 0 $X=7490 $Y=3230
X17 3 M2_M1_CDNS_7650569203814 $T=10320 3640 0 0 $X=10190 $Y=3510
X18 4 M2_M1_CDNS_7650569203815 $T=3420 5920 0 0 $X=3290 $Y=5790
X19 1 4 12 5 10 2 8 xor $T=4170 3810 0 0 $X=1950 $Y=1250
X20 10 4 9 5 6 3 8 xor $T=8070 3810 0 0 $X=5850 $Y=1250
X21 3 M3_M2_CDNS_7650569203821 $T=7300 3360 0 0 $X=7170 $Y=3230
X22 3 M3_M2_CDNS_7650569203821 $T=10110 3640 0 0 $X=9980 $Y=3510
X23 11 10 3 4 5 9 2 8 13 14
+ 15 16 fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 12 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 4 1 12 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 2 1 10 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 9 10 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 4 10 9 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 3 10 6 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 7 11 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 4 11 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mult_auto                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mult_auto 20 19 2 1 21 22 23 24 4 25
+ 32 78 103 108 114 115 116 117
** N=209 EP=18 FDC=576
X0 1 M4_M3_CDNS_765056920380 $T=530 48380 0 0 $X=170 $Y=47890
X1 2 M4_M3_CDNS_765056920380 $T=630 57160 0 0 $X=270 $Y=56670
X2 3 M2_M1_CDNS_765056920381 $T=6850 68930 0 0 $X=6770 $Y=68800
X3 4 M2_M1_CDNS_765056920381 $T=6860 78720 0 0 $X=6780 $Y=78590
X4 5 M2_M1_CDNS_765056920381 $T=7150 48200 0 0 $X=7070 $Y=48070
X5 6 M2_M1_CDNS_765056920381 $T=7150 57670 0 0 $X=7070 $Y=57540
X6 7 M2_M1_CDNS_765056920381 $T=15370 42570 0 0 $X=15290 $Y=42440
X7 8 M2_M1_CDNS_765056920381 $T=15470 62060 0 0 $X=15390 $Y=61930
X8 9 M2_M1_CDNS_765056920381 $T=15470 71890 0 0 $X=15390 $Y=71760
X9 10 M2_M1_CDNS_765056920381 $T=15480 52820 0 0 $X=15400 $Y=52690
X10 11 M2_M1_CDNS_765056920381 $T=36990 34960 0 0 $X=36910 $Y=34830
X11 12 M2_M1_CDNS_765056920381 $T=37850 43590 0 0 $X=37770 $Y=43460
X12 13 M2_M1_CDNS_765056920381 $T=39090 51720 0 0 $X=39010 $Y=51590
X13 14 M2_M1_CDNS_765056920381 $T=40940 59910 0 0 $X=40860 $Y=59780
X14 15 M2_M1_CDNS_765056920381 $T=63420 25360 0 0 $X=63340 $Y=25230
X15 16 M2_M1_CDNS_765056920381 $T=63680 34640 0 0 $X=63600 $Y=34510
X16 17 M2_M1_CDNS_765056920381 $T=64220 42710 0 0 $X=64140 $Y=42580
X17 18 M2_M1_CDNS_765056920381 $T=65650 50790 0 0 $X=65570 $Y=50660
X18 19 M3_M2_CDNS_765056920382 $T=3540 68870 0 0 $X=3460 $Y=68460
X19 20 M3_M2_CDNS_765056920382 $T=3540 78670 0 0 $X=3460 $Y=78260
X20 1 M3_M2_CDNS_765056920382 $T=3840 48140 0 0 $X=3760 $Y=47730
X21 2 M3_M2_CDNS_765056920382 $T=3840 57600 0 0 $X=3760 $Y=57190
X22 21 M3_M2_CDNS_765056920382 $T=4840 68580 0 0 $X=4760 $Y=68170
X23 21 M3_M2_CDNS_765056920382 $T=4840 78370 0 0 $X=4760 $Y=77960
X24 21 M3_M2_CDNS_765056920382 $T=5140 47840 0 0 $X=5060 $Y=47430
X25 21 M3_M2_CDNS_765056920382 $T=5140 57310 0 0 $X=5060 $Y=56900
X26 1 M3_M2_CDNS_765056920382 $T=12060 42520 0 0 $X=11980 $Y=42110
X27 2 M3_M2_CDNS_765056920382 $T=12160 52760 0 0 $X=12080 $Y=52350
X28 19 M3_M2_CDNS_765056920382 $T=12160 62010 0 0 $X=12080 $Y=61600
X29 20 M3_M2_CDNS_765056920382 $T=12160 71820 0 0 $X=12080 $Y=71410
X30 22 M3_M2_CDNS_765056920382 $T=13360 42210 0 0 $X=13280 $Y=41800
X31 22 M3_M2_CDNS_765056920382 $T=13460 52460 0 0 $X=13380 $Y=52050
X32 22 M3_M2_CDNS_765056920382 $T=13460 61710 0 0 $X=13380 $Y=61300
X33 22 M3_M2_CDNS_765056920382 $T=13460 71540 0 0 $X=13380 $Y=71130
X34 1 M3_M2_CDNS_765056920382 $T=33680 34900 0 0 $X=33600 $Y=34490
X35 2 M3_M2_CDNS_765056920382 $T=34530 43540 0 0 $X=34450 $Y=43130
X36 23 M3_M2_CDNS_765056920382 $T=34980 34600 0 0 $X=34900 $Y=34190
X37 19 M3_M2_CDNS_765056920382 $T=35730 51660 0 0 $X=35650 $Y=51250
X38 23 M3_M2_CDNS_765056920382 $T=35830 43240 0 0 $X=35750 $Y=42830
X39 23 M3_M2_CDNS_765056920382 $T=37030 51360 0 0 $X=36950 $Y=50950
X40 20 M3_M2_CDNS_765056920382 $T=37620 59850 0 0 $X=37540 $Y=59440
X41 23 M3_M2_CDNS_765056920382 $T=38920 59550 0 0 $X=38840 $Y=59140
X42 1 M3_M2_CDNS_765056920382 $T=60120 25320 0 0 $X=60040 $Y=24910
X43 2 M3_M2_CDNS_765056920382 $T=60360 34570 0 0 $X=60280 $Y=34160
X44 19 M3_M2_CDNS_765056920382 $T=60910 42670 0 0 $X=60830 $Y=42260
X45 24 M3_M2_CDNS_765056920382 $T=61420 25010 0 0 $X=61340 $Y=24600
X46 24 M3_M2_CDNS_765056920382 $T=61660 34270 0 0 $X=61580 $Y=33860
X47 24 M3_M2_CDNS_765056920382 $T=62210 42370 0 0 $X=62130 $Y=41960
X48 20 M3_M2_CDNS_765056920382 $T=62340 50730 0 0 $X=62260 $Y=50320
X49 24 M3_M2_CDNS_765056920382 $T=63640 50430 0 0 $X=63560 $Y=50020
X50 19 M2_M1_CDNS_765056920383 $T=3540 68870 0 0 $X=3460 $Y=68460
X51 20 M2_M1_CDNS_765056920383 $T=3540 78670 0 0 $X=3460 $Y=78260
X52 1 M2_M1_CDNS_765056920383 $T=3840 48140 0 0 $X=3760 $Y=47730
X53 2 M2_M1_CDNS_765056920383 $T=3840 57600 0 0 $X=3760 $Y=57190
X54 21 M2_M1_CDNS_765056920383 $T=4840 68580 0 0 $X=4760 $Y=68170
X55 21 M2_M1_CDNS_765056920383 $T=4840 78370 0 0 $X=4760 $Y=77960
X56 21 M2_M1_CDNS_765056920383 $T=5140 47840 0 0 $X=5060 $Y=47430
X57 21 M2_M1_CDNS_765056920383 $T=5140 57310 0 0 $X=5060 $Y=56900
X58 1 M2_M1_CDNS_765056920383 $T=12060 42520 0 0 $X=11980 $Y=42110
X59 2 M2_M1_CDNS_765056920383 $T=12160 52760 0 0 $X=12080 $Y=52350
X60 19 M2_M1_CDNS_765056920383 $T=12160 62010 0 0 $X=12080 $Y=61600
X61 20 M2_M1_CDNS_765056920383 $T=12160 71820 0 0 $X=12080 $Y=71410
X62 22 M2_M1_CDNS_765056920383 $T=13360 42210 0 0 $X=13280 $Y=41800
X63 22 M2_M1_CDNS_765056920383 $T=13460 52460 0 0 $X=13380 $Y=52050
X64 22 M2_M1_CDNS_765056920383 $T=13460 61710 0 0 $X=13380 $Y=61300
X65 22 M2_M1_CDNS_765056920383 $T=13460 71540 0 0 $X=13380 $Y=71130
X66 1 M2_M1_CDNS_765056920383 $T=33680 34900 0 0 $X=33600 $Y=34490
X67 2 M2_M1_CDNS_765056920383 $T=34530 43540 0 0 $X=34450 $Y=43130
X68 23 M2_M1_CDNS_765056920383 $T=34980 34600 0 0 $X=34900 $Y=34190
X69 19 M2_M1_CDNS_765056920383 $T=35730 51660 0 0 $X=35650 $Y=51250
X70 23 M2_M1_CDNS_765056920383 $T=35830 43240 0 0 $X=35750 $Y=42830
X71 23 M2_M1_CDNS_765056920383 $T=37030 51360 0 0 $X=36950 $Y=50950
X72 20 M2_M1_CDNS_765056920383 $T=37620 59850 0 0 $X=37540 $Y=59440
X73 23 M2_M1_CDNS_765056920383 $T=38920 59550 0 0 $X=38840 $Y=59140
X74 1 M2_M1_CDNS_765056920383 $T=60120 25320 0 0 $X=60040 $Y=24910
X75 2 M2_M1_CDNS_765056920383 $T=60360 34570 0 0 $X=60280 $Y=34160
X76 19 M2_M1_CDNS_765056920383 $T=60910 42670 0 0 $X=60830 $Y=42260
X77 24 M2_M1_CDNS_765056920383 $T=61420 25010 0 0 $X=61340 $Y=24600
X78 24 M2_M1_CDNS_765056920383 $T=61660 34270 0 0 $X=61580 $Y=33860
X79 24 M2_M1_CDNS_765056920383 $T=62210 42370 0 0 $X=62130 $Y=41960
X80 20 M2_M1_CDNS_765056920383 $T=62340 50730 0 0 $X=62260 $Y=50320
X81 24 M2_M1_CDNS_765056920383 $T=63640 50430 0 0 $X=63560 $Y=50020
X82 19 M4_M3_CDNS_765056920384 $T=550 69610 0 0 $X=110 $Y=69200
X83 20 M4_M3_CDNS_765056920384 $T=740 78860 0 0 $X=300 $Y=78450
X84 19 M4_M3_CDNS_765056920385 $T=3540 68870 0 0 $X=3460 $Y=68460
X85 20 M4_M3_CDNS_765056920385 $T=3540 78670 0 0 $X=3460 $Y=78260
X86 1 M4_M3_CDNS_765056920385 $T=3840 48140 0 0 $X=3760 $Y=47730
X87 2 M4_M3_CDNS_765056920385 $T=3840 57600 0 0 $X=3760 $Y=57190
X88 1 M4_M3_CDNS_765056920385 $T=12060 42520 0 0 $X=11980 $Y=42110
X89 20 M4_M3_CDNS_765056920385 $T=12150 71810 0 0 $X=12070 $Y=71400
X90 2 M4_M3_CDNS_765056920385 $T=12160 52760 0 0 $X=12080 $Y=52350
X91 19 M4_M3_CDNS_765056920385 $T=12160 62010 0 0 $X=12080 $Y=61600
X92 1 M4_M3_CDNS_765056920385 $T=33680 34900 0 0 $X=33600 $Y=34490
X93 2 M4_M3_CDNS_765056920385 $T=34530 43540 0 0 $X=34450 $Y=43130
X94 19 M4_M3_CDNS_765056920385 $T=35730 51660 0 0 $X=35650 $Y=51250
X95 20 M4_M3_CDNS_765056920385 $T=37620 59850 0 0 $X=37540 $Y=59440
X96 1 M4_M3_CDNS_765056920385 $T=60120 25320 0 0 $X=60040 $Y=24910
X97 2 M4_M3_CDNS_765056920385 $T=60360 34570 0 0 $X=60280 $Y=34160
X98 19 M4_M3_CDNS_765056920385 $T=60910 42670 0 0 $X=60830 $Y=42260
X99 20 M4_M3_CDNS_765056920385 $T=62340 50730 0 0 $X=62260 $Y=50320
X100 1 M5_M4_CDNS_765056920386 $T=33830 48370 0 0 $X=33750 $Y=48240
X101 2 M5_M4_CDNS_765056920386 $T=34690 57170 0 0 $X=34610 $Y=57040
X102 1 M5_M4_CDNS_765056920386 $T=35210 48370 0 0 $X=35130 $Y=48240
X103 19 M5_M4_CDNS_765056920386 $T=36060 69610 0 0 $X=35980 $Y=69480
X104 2 M5_M4_CDNS_765056920386 $T=36620 57170 0 0 $X=36540 $Y=57040
X105 19 M5_M4_CDNS_765056920386 $T=39250 69610 0 0 $X=39170 $Y=69480
X106 25 M5_M4_CDNS_765056920386 $T=59850 67350 0 0 $X=59770 $Y=67220
X107 25 M5_M4_CDNS_765056920386 $T=64530 67360 0 0 $X=64450 $Y=67230
X108 26 M4_M3_CDNS_765056920387 $T=34420 41500 0 0 $X=34340 $Y=41370
X109 27 M4_M3_CDNS_765056920387 $T=35180 50790 0 0 $X=35100 $Y=50660
X110 28 M4_M3_CDNS_765056920387 $T=36700 58320 0 0 $X=36620 $Y=58190
X111 25 M4_M3_CDNS_765056920387 $T=38150 67350 0 0 $X=38070 $Y=67220
X112 26 M4_M3_CDNS_765056920387 $T=39220 41500 0 0 $X=39140 $Y=41370
X113 27 M4_M3_CDNS_765056920387 $T=40000 50780 0 0 $X=39920 $Y=50650
X114 28 M4_M3_CDNS_765056920387 $T=43090 58320 0 0 $X=43010 $Y=58190
X115 29 M4_M3_CDNS_765056920387 $T=60680 32400 0 0 $X=60600 $Y=32270
X116 30 M4_M3_CDNS_765056920387 $T=60890 40780 0 0 $X=60810 $Y=40650
X117 31 M4_M3_CDNS_765056920387 $T=61780 49010 0 0 $X=61700 $Y=48880
X118 32 M4_M3_CDNS_765056920387 $T=62920 58800 0 0 $X=62840 $Y=58670
X119 29 M4_M3_CDNS_765056920387 $T=65120 32400 0 0 $X=65040 $Y=32270
X120 30 M4_M3_CDNS_765056920387 $T=66260 40780 0 0 $X=66180 $Y=40650
X121 31 M4_M3_CDNS_765056920387 $T=67200 49000 0 0 $X=67120 $Y=48870
X122 32 M4_M3_CDNS_765056920387 $T=86280 63220 0 0 $X=86200 $Y=63090
X123 25 M4_M3_CDNS_765056920387 $T=87220 73220 0 0 $X=87140 $Y=73090
X124 7 M3_M2_CDNS_765056920388 $T=15370 42570 0 0 $X=15290 $Y=42440
X125 10 M3_M2_CDNS_765056920388 $T=19170 51720 0 0 $X=19090 $Y=51590
X126 5 M3_M2_CDNS_765056920388 $T=19210 50780 0 0 $X=19130 $Y=50650
X127 6 M3_M2_CDNS_765056920388 $T=20100 59120 0 0 $X=20020 $Y=58990
X128 8 M3_M2_CDNS_765056920388 $T=20110 60060 0 0 $X=20030 $Y=59930
X129 9 M3_M2_CDNS_765056920388 $T=22540 68220 0 0 $X=22460 $Y=68090
X130 3 M3_M2_CDNS_765056920388 $T=22550 67750 0 0 $X=22470 $Y=67620
X131 12 M3_M2_CDNS_765056920388 $T=39390 43590 0 0 $X=39310 $Y=43460
X132 11 M3_M2_CDNS_765056920388 $T=39400 34950 0 0 $X=39320 $Y=34820
X133 13 M3_M2_CDNS_765056920388 $T=41300 51720 0 0 $X=41220 $Y=51590
X134 14 M3_M2_CDNS_765056920388 $T=43140 59910 0 0 $X=43060 $Y=59780
X135 16 M3_M2_CDNS_765056920388 $T=66170 34680 0 0 $X=66090 $Y=34550
X136 15 M3_M2_CDNS_765056920388 $T=66360 26140 0 0 $X=66280 $Y=26010
X137 17 M3_M2_CDNS_765056920388 $T=66510 43080 0 0 $X=66430 $Y=42950
X138 18 M3_M2_CDNS_765056920388 $T=68160 51630 0 0 $X=68080 $Y=51500
X139 19 33 21 34 3 35 174 118 and2 $T=5890 68510 0 0 $X=3220 $Y=65930
X140 20 36 21 37 4 35 175 119 and2 $T=5890 78310 0 0 $X=3220 $Y=75730
X141 1 38 21 39 5 35 176 120 and2 $T=6190 47780 0 0 $X=3520 $Y=45200
X142 2 40 21 41 6 35 177 121 and2 $T=6190 57250 0 0 $X=3520 $Y=54670
X143 1 42 22 43 7 35 178 122 and2 $T=14410 42150 0 0 $X=11740 $Y=39570
X144 2 44 22 45 10 35 179 123 and2 $T=14510 52400 0 0 $X=11840 $Y=49820
X145 19 46 22 47 8 35 180 124 and2 $T=14510 61650 0 0 $X=11840 $Y=59070
X146 20 48 22 49 9 35 181 125 and2 $T=14510 71470 0 0 $X=11840 $Y=68890
X147 1 50 23 51 11 35 182 126 and2 $T=36030 34540 0 0 $X=33360 $Y=31960
X148 2 52 23 53 12 35 183 127 and2 $T=36880 43180 0 0 $X=34210 $Y=40600
X149 19 54 23 55 13 35 184 128 and2 $T=38080 51300 0 0 $X=35410 $Y=48720
X150 20 56 23 57 14 35 185 129 and2 $T=39970 59490 0 0 $X=37300 $Y=56910
X151 1 58 24 59 15 35 186 130 and2 $T=62470 24950 0 0 $X=59800 $Y=22370
X152 2 60 24 61 16 35 187 131 and2 $T=62710 34210 0 0 $X=60040 $Y=31630
X153 19 62 24 63 17 35 188 132 and2 $T=63260 42310 0 0 $X=60590 $Y=39730
X154 20 64 24 65 18 35 189 133 and2 $T=64690 50370 0 0 $X=62020 $Y=47790
X155 66 7 67 68 26 69 35 134 half_adder $T=19950 40210 0 0 $X=22250 $Y=40490
X156 9 3 70 71 25 72 35 136 half_adder $T=20250 64650 0 0 $X=22550 $Y=64930
X157 14 28 73 74 32 75 35 138 half_adder $T=45360 56090 0 0 $X=47660 $Y=56370
X158 18 31 76 77 78 79 35 140 half_adder $T=69570 48090 0 0 $X=71870 $Y=48370
X159 10 5 80 81 35 27 82 35 144 143
+ 145 142 full_adder $T=18880 47880 0 0 $X=20660 $Y=49130
X160 8 6 83 84 85 28 86 35 148 147
+ 149 146 full_adder $T=18880 56220 0 0 $X=20660 $Y=57470
X161 12 26 87 88 89 30 90 35 152 151
+ 153 150 full_adder $T=43990 39660 0 0 $X=45770 $Y=40910
X162 13 27 91 92 93 31 94 35 156 155
+ 157 154 full_adder $T=43990 47880 0 0 $X=45770 $Y=49130
X163 11 95 96 97 98 29 99 35 160 159
+ 161 158 full_adder $T=44590 31440 0 0 $X=46370 $Y=32690
X164 17 30 100 101 102 103 104 35 164 163
+ 165 162 full_adder $T=69190 39320 0 0 $X=70970 $Y=40570
X165 16 29 105 106 107 108 109 35 168 167
+ 169 166 full_adder $T=69850 30860 0 0 $X=71630 $Y=32110
X166 15 110 111 112 113 114 115 35 172 171
+ 173 170 full_adder $T=69860 22410 0 0 $X=71640 $Y=23660
M0 118 19 33 33 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3640 $Y=69440 $dt=1
M1 119 20 36 36 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3640 $Y=79240 $dt=1
M2 120 1 38 38 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3940 $Y=48710 $dt=1
M3 121 2 40 40 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3940 $Y=58180 $dt=1
M4 33 19 118 33 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4050 $Y=69440 $dt=1
M5 36 20 119 36 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4050 $Y=79240 $dt=1
M6 38 1 120 38 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4350 $Y=48710 $dt=1
M7 40 2 121 40 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4350 $Y=58180 $dt=1
M8 118 21 33 33 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4940 $Y=69440 $dt=1
M9 119 21 36 36 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4940 $Y=79240 $dt=1
M10 120 21 38 38 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=5240 $Y=48710 $dt=1
M11 121 21 40 40 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=5240 $Y=58180 $dt=1
M12 122 1 42 42 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12160 $Y=43080 $dt=1
M13 123 2 44 44 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=53330 $dt=1
M14 124 19 46 46 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=62580 $dt=1
M15 125 20 48 48 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=72400 $dt=1
M16 42 1 122 42 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12570 $Y=43080 $dt=1
M17 44 2 123 44 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=53330 $dt=1
M18 46 19 124 46 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=62580 $dt=1
M19 48 20 125 48 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=72400 $dt=1
M20 122 22 42 42 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13460 $Y=43080 $dt=1
M21 123 22 44 44 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=53330 $dt=1
M22 124 22 46 46 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=62580 $dt=1
M23 125 22 48 48 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=72400 $dt=1
M24 126 1 50 50 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=33780 $Y=35470 $dt=1
M25 50 1 126 50 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=34190 $Y=35470 $dt=1
M26 127 2 52 52 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=34630 $Y=44110 $dt=1
M27 52 2 127 52 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=35040 $Y=44110 $dt=1
M28 126 23 50 50 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=35080 $Y=35470 $dt=1
M29 128 19 54 54 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=35830 $Y=52230 $dt=1
M30 127 23 52 52 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=35930 $Y=44110 $dt=1
M31 54 19 128 54 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=36240 $Y=52230 $dt=1
M32 128 23 54 54 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=37130 $Y=52230 $dt=1
M33 129 20 56 56 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=37720 $Y=60420 $dt=1
M34 56 20 129 56 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=38130 $Y=60420 $dt=1
M35 129 23 56 56 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=39020 $Y=60420 $dt=1
M36 130 1 58 58 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=60220 $Y=25880 $dt=1
M37 131 2 60 60 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=60460 $Y=35140 $dt=1
M38 58 1 130 58 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=60630 $Y=25880 $dt=1
M39 60 2 131 60 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=60870 $Y=35140 $dt=1
M40 132 19 62 62 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=61010 $Y=43240 $dt=1
M41 62 19 132 62 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=61420 $Y=43240 $dt=1
M42 130 24 58 58 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=61520 $Y=25880 $dt=1
M43 131 24 60 60 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=61760 $Y=35140 $dt=1
M44 132 24 62 62 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=62310 $Y=43240 $dt=1
M45 133 20 64 64 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=62440 $Y=51300 $dt=1
M46 64 20 133 64 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=62850 $Y=51300 $dt=1
M47 133 24 64 64 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=63740 $Y=51300 $dt=1
.ends mult_auto
