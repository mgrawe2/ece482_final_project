* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : half_adder                                   *
* Netlisted  : Sat Dec  6 11:38:36 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765042711150                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765042711150 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765042711150

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765042711151                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765042711151 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765042711151

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765042711152                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765042711152 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765042711152

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765042711153                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765042711153 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765042711153

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_765042711154                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_765042711154 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_765042711154

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765042711155                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765042711155 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765042711155

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_765042711156                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_765042711156 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_765042711156

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765042711157                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765042711157 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765042711157

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765042711150                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765042711150 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765042711150

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765042711151                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765042711151 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_765042711151

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765042711152                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765042711152 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765042711152

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X0 3 M1_NWELL_CDNS_765042711154 $T=190 2570 0 0 $X=-230 $Y=2270
X1 4 M1_PSUB_CDNS_765042711156 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 1 M1_PO_CDNS_765042711157 $T=-160 30 0 0 $X=-260 $Y=-330
X3 3 2 1 3 4 3 pmos1v_CDNS_765042711151 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 2 1 4 4 nmos1v_CDNS_765042711152 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7
** N=7 EP=7 FDC=12
X0 1 M1_NWELL_CDNS_765042711154 $T=-1350 2870 0 0 $X=-1770 $Y=2570
X1 6 M2_M1_CDNS_765042711155 $T=-2410 -1220 0 0 $X=-2490 $Y=-1470
X2 7 M2_M1_CDNS_765042711155 $T=-2000 1650 0 0 $X=-2080 $Y=1400
X3 6 M2_M1_CDNS_765042711155 $T=-1590 -1220 0 0 $X=-1670 $Y=-1470
X4 6 M2_M1_CDNS_765042711155 $T=-1110 -1220 0 0 $X=-1190 $Y=-1470
X5 7 M2_M1_CDNS_765042711155 $T=-700 1650 0 0 $X=-780 $Y=1400
X6 6 M2_M1_CDNS_765042711155 $T=-290 -1220 0 0 $X=-370 $Y=-1470
X7 4 M1_PSUB_CDNS_765042711156 $T=-700 -2440 0 0 $X=-1080 $Y=-2580
X8 2 M1_PO_CDNS_765042711157 $T=-2350 360 0 0 $X=-2450 $Y=0
X9 3 M1_PO_CDNS_765042711157 $T=-1050 60 0 0 $X=-1150 $Y=-300
X10 6 6 7 2 4 nmos1v_CDNS_765042711150 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 6 6 4 3 4 nmos1v_CDNS_765042711150 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X12 1 7 2 1 4 1 pmos1v_CDNS_765042711151 $T=-2250 930 0 0 $X=-2670 $Y=730
X13 1 7 3 1 4 1 pmos1v_CDNS_765042711151 $T=-950 930 0 0 $X=-1370 $Y=730
X14 7 5 1 4 inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 7 2 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-2250 $Y=930 $dt=1
M1 1 2 7 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-1840 $Y=930 $dt=1
M2 7 3 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-950 $Y=930 $dt=1
M3 1 3 7 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M4 5 7 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M5 1 7 5 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7650427111510                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7650427111510 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7650427111510

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
** N=6 EP=6 FDC=12
X0 5 M2_M1_CDNS_765042711150 $T=-30 -450 0 0 $X=-160 $Y=-580
X1 6 M2_M1_CDNS_765042711150 $T=1330 -190 0 0 $X=1200 $Y=-320
X2 5 M2_M1_CDNS_765042711151 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X3 5 M2_M1_CDNS_765042711151 $T=-250 380 0 0 $X=-380 $Y=250
X4 6 M2_M1_CDNS_765042711155 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X5 6 M2_M1_CDNS_765042711155 $T=-660 950 0 0 $X=-740 $Y=700
X6 6 M2_M1_CDNS_765042711155 $T=160 -1560 0 0 $X=80 $Y=-1810
X7 6 M2_M1_CDNS_765042711155 $T=160 950 0 0 $X=80 $Y=700
X8 6 M2_M1_CDNS_765042711155 $T=1050 -1560 0 0 $X=970 $Y=-1810
X9 6 M2_M1_CDNS_765042711155 $T=1050 950 0 0 $X=970 $Y=700
X10 6 5 1 6 3 4 pmos1v_CDNS_765042711151 $T=-500 230 0 0 $X=-920 $Y=30
X11 1 6 5 1 3 4 pmos1v_CDNS_765042711151 $T=800 230 0 0 $X=380 $Y=30
X12 6 5 2 6 3 nmos1v_CDNS_765042711152 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X13 2 6 5 2 3 nmos1v_CDNS_765042711152 $T=800 -1920 0 0 $X=380 $Y=-2120
X14 1 2 4 3 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
X15 1 M1_PO_CDNS_7650427111510 $T=-450 10 0 0 $X=-550 $Y=-110
X16 1 M1_PO_CDNS_7650427111510 $T=-450 1890 0 0 $X=-550 $Y=1770
X17 2 M1_PO_CDNS_7650427111510 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X18 1 M1_PO_CDNS_7650427111510 $T=-40 1890 0 0 $X=-140 $Y=1770
X19 5 M1_PO_CDNS_7650427111510 $T=850 -980 0 0 $X=750 $Y=-1100
M0 2 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1800 $Y=230 $dt=1
M1 4 1 2 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1390 $Y=230 $dt=1
M2 5 1 6 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-500 $Y=230 $dt=1
M3 6 1 5 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M4 6 5 1 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M5 1 5 6 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 3 1 4 2 5 6
** N=9 EP=6 FDC=24
X0 1 M2_M1_CDNS_765042711150 $T=2760 2580 0 0 $X=2630 $Y=2450
X1 1 M2_M1_CDNS_765042711150 $T=7960 2810 0 0 $X=7830 $Y=2680
X2 2 M2_M1_CDNS_765042711151 $T=6360 3430 0 0 $X=6230 $Y=3300
X3 1 M3_M2_CDNS_765042711152 $T=2760 3570 0 0 $X=2680 $Y=3440
X4 3 M3_M2_CDNS_765042711152 $T=4630 3110 0 0 $X=4550 $Y=2980
X5 4 M3_M2_CDNS_765042711152 $T=9970 3310 0 0 $X=9890 $Y=3180
X6 2 M3_M2_CDNS_765042711152 $T=10180 2730 0 0 $X=10100 $Y=2600
X7 4 M2_M1_CDNS_765042711153 $T=9970 3310 0 0 $X=9890 $Y=3180
X8 2 M2_M1_CDNS_765042711153 $T=10180 2730 0 0 $X=10100 $Y=2600
X9 5 3 1 6 4 9 8 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X10 1 7 6 5 3 2 xor $T=4660 3560 0 0 $X=2440 $Y=1000
.ends half_adder
