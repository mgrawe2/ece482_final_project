* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : and2                                         *
* Netlisted  : Thu Dec  4 17:31:13 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764891067850                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764891067850 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764891067850

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764891067851                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764891067851 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764891067851

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764891067852                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764891067852 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_764891067852

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764891067853                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764891067853 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764891067853

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_764891067854                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_764891067854 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_764891067854

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764891067855                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764891067855 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764891067855

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764891067850                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764891067850 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764891067850

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764891067851                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764891067851 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_764891067851

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand2                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand2 1 2 3 4 5 6
** N=6 EP=6 FDC=8
X0 3 M1_NWELL_CDNS_764891067852 $T=1290 2080 0 0 $X=870 $Y=1780
X1 6 M2_M1_CDNS_764891067853 $T=230 -2010 0 0 $X=150 $Y=-2260
X2 1 M2_M1_CDNS_764891067853 $T=640 860 0 0 $X=560 $Y=610
X3 6 M2_M1_CDNS_764891067853 $T=1050 -2010 0 0 $X=970 $Y=-2260
X4 6 M2_M1_CDNS_764891067853 $T=1530 -2010 0 0 $X=1450 $Y=-2260
X5 1 M2_M1_CDNS_764891067853 $T=1940 860 0 0 $X=1860 $Y=610
X6 6 M2_M1_CDNS_764891067853 $T=2350 -2010 0 0 $X=2270 $Y=-2260
X7 5 M1_PSUB_CDNS_764891067854 $T=1940 -3230 0 0 $X=1560 $Y=-3370
X8 2 M1_PO_CDNS_764891067855 $T=290 -430 0 0 $X=190 $Y=-790
X9 4 M1_PO_CDNS_764891067855 $T=1590 -730 0 0 $X=1490 $Y=-1090
X10 6 6 1 2 5 nmos1v_CDNS_764891067850 $T=390 -2730 0 0 $X=-30 $Y=-2930
X11 6 6 5 4 5 nmos1v_CDNS_764891067850 $T=1690 -2730 0 0 $X=1270 $Y=-2930
X12 1 3 3 2 5 3 pmos1v_CDNS_764891067851 $T=390 140 0 0 $X=-30 $Y=-60
X13 1 3 3 4 5 3 pmos1v_CDNS_764891067851 $T=1690 140 0 0 $X=1270 $Y=-60
M0 1 2 3 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=390 $Y=140 $dt=1
M1 3 2 1 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=800 $Y=140 $dt=1
M2 1 4 3 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1690 $Y=140 $dt=1
M3 3 4 1 3 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=2100 $Y=140 $dt=1
.ends nand2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764891067852                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764891067852 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 4 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 3 4 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764891067852

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
** N=4 EP=4 FDC=4
X0 1 M1_NWELL_CDNS_764891067852 $T=190 2570 0 0 $X=-230 $Y=2270
X1 2 M1_PSUB_CDNS_764891067854 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 3 M1_PO_CDNS_764891067855 $T=-160 30 0 0 $X=-260 $Y=-330
X3 4 1 1 3 2 1 pmos1v_CDNS_764891067851 $T=-60 630 0 0 $X=-480 $Y=430
X4 2 4 2 3 2 nmos1v_CDNS_764891067852 $T=-60 -1520 0 0 $X=-480 $Y=-1720
M0 4 3 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-60 $Y=630 $dt=1
M1 1 3 4 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=350 $Y=630 $dt=1
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 5 6
** N=7 EP=5 FDC=12
X0 1 M2_M1_CDNS_764891067850 $T=-2340 370 0 0 $X=-2420 $Y=100
X1 2 M2_M1_CDNS_764891067850 $T=-1050 50 0 0 $X=-1130 $Y=-220
X2 3 M2_M1_CDNS_764891067850 $T=1110 410 0 0 $X=1030 $Y=140
X3 1 M3_M2_CDNS_764891067851 $T=-2340 370 0 0 $X=-2420 $Y=100
X4 2 M3_M2_CDNS_764891067851 $T=-1050 50 0 0 $X=-1130 $Y=-220
X5 3 M3_M2_CDNS_764891067851 $T=1110 410 0 0 $X=1030 $Y=140
X6 4 1 5 2 6 7 nand2 $T=-2640 790 0 0 $X=-2670 $Y=-2580
X7 5 6 4 3 inv $T=410 300 0 0 $X=-70 $Y=-1860
.ends and2
