* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mult_auto                                    *
* Netlisted  : Sat Dec  6 18:47:50 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765068464210                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765068464210 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765068464210

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765068464211                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765068464211 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765068464211

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765068464212                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765068464212 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765068464212

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765068464213                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765068464213 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765068464213

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765068464214                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765068464214 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765068464214

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765068464215                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765068464215 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765068464215

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765068464216                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765068464216 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765068464216

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765068464217                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765068464217 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765068464217

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765068464218                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765068464218 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765068464218

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765068464219                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765068464219 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765068464219

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7650684642110                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7650684642110 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7650684642110

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7650684642111                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7650684642111 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7650684642111

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7650684642113                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7650684642113 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7650684642113

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7650684642114                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7650684642114 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7650684642114

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7650684642115                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7650684642115 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7650684642115

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_7650684642116                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_7650684642116 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_7650684642116

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_7650684642117                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_7650684642117 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_7650684642117

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_7650684642118                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_7650684642118 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_7650684642118

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_7650684642119                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_7650684642119 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_7650684642119

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_7650684642120                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_7650684642120 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_7650684642120

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7650684642121                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7650684642121 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7650684642121

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_7650684642122                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_7650684642122 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_7650684642122

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7650684642123                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7650684642123 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7650684642123

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765068464210                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765068464210 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765068464210

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765068464211                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765068464211 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_765068464211

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765068464212                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765068464212 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765068464212

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X0 2 M1_NWELL_CDNS_7650684642120 $T=190 2570 0 0 $X=-230 $Y=2270
X1 4 M1_PSUB_CDNS_7650684642122 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 1 M1_PO_CDNS_7650684642123 $T=-160 30 0 0 $X=-260 $Y=-330
X3 2 3 1 2 4 2 pmos1v_CDNS_765068464211 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 3 1 4 4 nmos1v_CDNS_765068464212 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=9
X0 2 M1_NWELL_CDNS_7650684642120 $T=-1350 2870 0 0 $X=-1770 $Y=2570
X1 6 M2_M1_CDNS_7650684642121 $T=-2410 -1220 0 0 $X=-2490 $Y=-1470
X2 7 M2_M1_CDNS_7650684642121 $T=-2000 1650 0 0 $X=-2080 $Y=1400
X3 6 M2_M1_CDNS_7650684642121 $T=-1590 -1220 0 0 $X=-1670 $Y=-1470
X4 6 M2_M1_CDNS_7650684642121 $T=-1110 -1220 0 0 $X=-1190 $Y=-1470
X5 7 M2_M1_CDNS_7650684642121 $T=-700 1650 0 0 $X=-780 $Y=1400
X6 6 M2_M1_CDNS_7650684642121 $T=-290 -1220 0 0 $X=-370 $Y=-1470
X7 4 M1_PSUB_CDNS_7650684642122 $T=-700 -2440 0 0 $X=-1080 $Y=-2580
X8 1 M1_PO_CDNS_7650684642123 $T=-2350 360 0 0 $X=-2450 $Y=0
X9 3 M1_PO_CDNS_7650684642123 $T=-1050 60 0 0 $X=-1150 $Y=-300
X10 6 6 7 1 4 nmos1v_CDNS_765068464210 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 6 6 4 3 4 nmos1v_CDNS_765068464210 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X12 2 7 1 2 4 2 pmos1v_CDNS_765068464211 $T=-2250 930 0 0 $X=-2670 $Y=730
X13 2 7 3 2 4 2 pmos1v_CDNS_765068464211 $T=-950 930 0 0 $X=-1370 $Y=730
X14 7 2 5 4 inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 2 3 7 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M1 5 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M2 2 7 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7650684642124                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7650684642124 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7650684642124

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7650684642125                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7650684642125 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7650684642125

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7650684642128                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7650684642128 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7650684642128

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X0 5 M2_M1_CDNS_7650684642121 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X1 5 M2_M1_CDNS_7650684642121 $T=-660 950 0 0 $X=-740 $Y=700
X2 5 M2_M1_CDNS_7650684642121 $T=160 -1560 0 0 $X=80 $Y=-1810
X3 5 M2_M1_CDNS_7650684642121 $T=160 950 0 0 $X=80 $Y=700
X4 5 M2_M1_CDNS_7650684642121 $T=1050 -1560 0 0 $X=970 $Y=-1810
X5 5 M2_M1_CDNS_7650684642121 $T=1050 950 0 0 $X=970 $Y=700
X6 5 6 1 5 3 2 pmos1v_CDNS_765068464211 $T=-500 230 0 0 $X=-920 $Y=30
X7 1 5 6 1 3 2 pmos1v_CDNS_765068464211 $T=800 230 0 0 $X=380 $Y=30
X8 5 6 4 5 3 nmos1v_CDNS_765068464212 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X9 4 5 6 4 3 nmos1v_CDNS_765068464212 $T=800 -1920 0 0 $X=380 $Y=-2120
X10 1 2 4 3 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
X11 6 M2_M1_CDNS_7650684642124 $T=-30 -450 0 0 $X=-160 $Y=-580
X12 5 M2_M1_CDNS_7650684642124 $T=1330 -190 0 0 $X=1200 $Y=-320
X13 6 M2_M1_CDNS_7650684642125 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X14 6 M2_M1_CDNS_7650684642125 $T=-250 380 0 0 $X=-380 $Y=250
X15 1 M1_PO_CDNS_7650684642128 $T=-450 10 0 0 $X=-550 $Y=-110
X16 1 M1_PO_CDNS_7650684642128 $T=-450 1890 0 0 $X=-550 $Y=1770
X17 4 M1_PO_CDNS_7650684642128 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X18 1 M1_PO_CDNS_7650684642128 $T=-40 1890 0 0 $X=-140 $Y=1770
X19 6 M1_PO_CDNS_7650684642128 $T=850 -980 0 0 $X=750 $Y=-1100
M0 5 1 6 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 5 6 1 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 1 6 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 7
** N=9 EP=7 FDC=24
X0 6 M2_M1_CDNS_765068464211 $T=9970 3310 0 0 $X=9890 $Y=3180
X1 5 M2_M1_CDNS_765068464211 $T=10180 2730 0 0 $X=10100 $Y=2600
X2 1 M3_M2_CDNS_7650684642111 $T=2760 3570 0 0 $X=2680 $Y=3440
X3 2 M3_M2_CDNS_7650684642111 $T=4630 3110 0 0 $X=4550 $Y=2980
X4 6 M3_M2_CDNS_7650684642111 $T=9970 3310 0 0 $X=9890 $Y=3180
X5 5 M3_M2_CDNS_7650684642111 $T=10180 2730 0 0 $X=10100 $Y=2600
X6 2 4 1 3 6 9 8 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X7 1 M2_M1_CDNS_7650684642124 $T=2760 2580 0 0 $X=2630 $Y=2450
X8 1 M2_M1_CDNS_7650684642124 $T=7960 2810 0 0 $X=7830 $Y=2680
X9 5 M2_M1_CDNS_7650684642125 $T=6360 3430 0 0 $X=6230 $Y=3300
X10 1 4 3 7 5 2 xor $T=4660 3560 0 0 $X=2440 $Y=1000
M0 7 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2860 $Y=3790 $dt=1
M1 4 1 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3270 $Y=3790 $dt=1
M2 2 1 5 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4160 $Y=3790 $dt=1
M3 8 2 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6760 $Y=3790 $dt=1
M4 4 2 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7170 $Y=3790 $dt=1
M5 8 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8060 $Y=3790 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7650684642131                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7650684642131 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7650684642131

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765068464213                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765068464213 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_765068464213

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765068464214                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765068464214 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_765068464214

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=8
X0 1 M2_M1_CDNS_765068464211 $T=-830 -970 0 0 $X=-910 $Y=-1100
X1 2 M2_M1_CDNS_765068464211 $T=-220 -60 0 0 $X=-300 $Y=-190
X2 2 M2_M1_CDNS_765068464211 $T=200 730 0 0 $X=120 $Y=600
X3 1 M2_M1_CDNS_765068464211 $T=810 -970 0 0 $X=730 $Y=-1100
X4 4 M1_NWELL_CDNS_7650684642120 $T=-10 2990 0 0 $X=-430 $Y=2690
X5 5 M1_PSUB_CDNS_7650684642122 $T=0 -1600 0 0 $X=-380 $Y=-1740
X6 3 M1_PO_CDNS_7650684642123 $T=-590 550 0 0 $X=-690 $Y=190
X7 7 M1_PO_CDNS_7650684642123 $T=570 550 0 0 $X=470 $Y=190
X8 2 M1_PO_CDNS_7650684642128 $T=-220 -60 0 0 $X=-320 $Y=-180
X9 6 M1_PO_CDNS_7650684642128 $T=-210 730 0 0 $X=-310 $Y=610
X10 6 M1_PO_CDNS_7650684642128 $T=190 -60 0 0 $X=90 $Y=-180
X11 2 M1_PO_CDNS_7650684642128 $T=200 730 0 0 $X=100 $Y=610
X12 1 8 3 5 9 2 6 1 7 nmos1v_CDNS_765068464213 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 1 10 4 3 6 11 1 2 7 5
+ 4 pmos1v_CDNS_765068464214 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 1 2 3 4 5 6 7 8 9 10
+ 11
** N=15 EP=11 FDC=36
X0 2 M2_M1_CDNS_765068464211 $T=5250 3070 0 0 $X=5170 $Y=2940
X1 8 M2_M1_CDNS_765068464211 $T=9530 2380 0 0 $X=9450 $Y=2250
X2 9 M2_M1_CDNS_765068464211 $T=9530 5090 0 0 $X=9450 $Y=4960
X3 4 M2_M1_CDNS_765068464211 $T=10820 5970 0 0 $X=10740 $Y=5840
X4 8 M2_M1_CDNS_765068464211 $T=11040 2940 0 0 $X=10960 $Y=2810
X5 2 M2_M1_CDNS_765068464211 $T=11390 3320 0 0 $X=11310 $Y=3190
X6 7 M2_M1_CDNS_765068464211 $T=12920 3510 0 0 $X=12840 $Y=3380
X7 2 M4_M3_CDNS_7650684642110 $T=6980 3080 0 0 $X=6900 $Y=2950
X8 2 M4_M3_CDNS_7650684642110 $T=10140 2970 0 0 $X=10060 $Y=2840
X9 1 M3_M2_CDNS_7650684642111 $T=2270 3860 0 0 $X=2190 $Y=3730
X10 2 M3_M2_CDNS_7650684642111 $T=5790 3080 0 0 $X=5710 $Y=2950
X11 6 M3_M2_CDNS_7650684642111 $T=9120 4760 0 0 $X=9040 $Y=4630
X12 2 M3_M2_CDNS_7650684642111 $T=11410 2940 0 0 $X=11330 $Y=2810
X13 7 M3_M2_CDNS_7650684642111 $T=12920 3510 0 0 $X=12840 $Y=3380
X14 10 4 7 5 inv $T=12350 3410 0 0 $X=11870 $Y=1250
X15 4 M2_M1_CDNS_7650684642124 $T=6470 5920 0 0 $X=6340 $Y=5790
X16 3 M2_M1_CDNS_7650684642124 $T=7620 3360 0 0 $X=7490 $Y=3230
X17 3 M2_M1_CDNS_7650684642124 $T=10320 3640 0 0 $X=10190 $Y=3510
X18 4 M2_M1_CDNS_7650684642125 $T=3420 5920 0 0 $X=3290 $Y=5790
X19 1 4 5 11 9 2 xor $T=4170 3810 0 0 $X=1950 $Y=1250
X20 9 4 5 8 6 3 xor $T=8070 3810 0 0 $X=5850 $Y=1250
X21 3 M3_M2_CDNS_7650684642131 $T=7300 3360 0 0 $X=7170 $Y=3230
X22 3 M3_M2_CDNS_7650684642131 $T=10110 3640 0 0 $X=9980 $Y=3510
X23 10 9 3 4 5 8 2 12 13 14
+ 15 fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 11 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 4 1 11 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 2 1 9 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 8 9 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 4 9 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 3 9 6 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 7 10 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 4 10 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mult_auto                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mult_auto 20 19 2 1 21 22 23 24 4 28
+ 35 47 48 49 50 51 26 25
** N=143 EP=18 FDC=576
X0 1 M4_M3_CDNS_765068464210 $T=530 48380 0 0 $X=170 $Y=47890
X1 2 M4_M3_CDNS_765068464210 $T=630 57160 0 0 $X=270 $Y=56670
X2 3 M2_M1_CDNS_765068464211 $T=6850 68930 0 0 $X=6770 $Y=68800
X3 4 M2_M1_CDNS_765068464211 $T=6860 78720 0 0 $X=6780 $Y=78590
X4 5 M2_M1_CDNS_765068464211 $T=7150 48200 0 0 $X=7070 $Y=48070
X5 6 M2_M1_CDNS_765068464211 $T=7150 57670 0 0 $X=7070 $Y=57540
X6 7 M2_M1_CDNS_765068464211 $T=15370 42570 0 0 $X=15290 $Y=42440
X7 8 M2_M1_CDNS_765068464211 $T=15470 62060 0 0 $X=15390 $Y=61930
X8 9 M2_M1_CDNS_765068464211 $T=15470 71890 0 0 $X=15390 $Y=71760
X9 10 M2_M1_CDNS_765068464211 $T=15480 52820 0 0 $X=15400 $Y=52690
X10 11 M2_M1_CDNS_765068464211 $T=36990 34960 0 0 $X=36910 $Y=34830
X11 12 M2_M1_CDNS_765068464211 $T=37850 43590 0 0 $X=37770 $Y=43460
X12 13 M2_M1_CDNS_765068464211 $T=39090 51720 0 0 $X=39010 $Y=51590
X13 14 M2_M1_CDNS_765068464211 $T=40940 59910 0 0 $X=40860 $Y=59780
X14 15 M2_M1_CDNS_765068464211 $T=63420 25360 0 0 $X=63340 $Y=25230
X15 16 M2_M1_CDNS_765068464211 $T=63680 34640 0 0 $X=63600 $Y=34510
X16 17 M2_M1_CDNS_765068464211 $T=64220 42710 0 0 $X=64140 $Y=42580
X17 18 M2_M1_CDNS_765068464211 $T=65650 50790 0 0 $X=65570 $Y=50660
X18 19 M3_M2_CDNS_765068464212 $T=3540 68870 0 0 $X=3460 $Y=68460
X19 20 M3_M2_CDNS_765068464212 $T=3540 78670 0 0 $X=3460 $Y=78260
X20 1 M3_M2_CDNS_765068464212 $T=3840 48140 0 0 $X=3760 $Y=47730
X21 2 M3_M2_CDNS_765068464212 $T=3840 57600 0 0 $X=3760 $Y=57190
X22 21 M3_M2_CDNS_765068464212 $T=4840 68580 0 0 $X=4760 $Y=68170
X23 21 M3_M2_CDNS_765068464212 $T=4840 78370 0 0 $X=4760 $Y=77960
X24 21 M3_M2_CDNS_765068464212 $T=5140 47840 0 0 $X=5060 $Y=47430
X25 21 M3_M2_CDNS_765068464212 $T=5140 57310 0 0 $X=5060 $Y=56900
X26 1 M3_M2_CDNS_765068464212 $T=12060 42520 0 0 $X=11980 $Y=42110
X27 2 M3_M2_CDNS_765068464212 $T=12160 52760 0 0 $X=12080 $Y=52350
X28 19 M3_M2_CDNS_765068464212 $T=12160 62010 0 0 $X=12080 $Y=61600
X29 20 M3_M2_CDNS_765068464212 $T=12160 71820 0 0 $X=12080 $Y=71410
X30 22 M3_M2_CDNS_765068464212 $T=13360 42210 0 0 $X=13280 $Y=41800
X31 22 M3_M2_CDNS_765068464212 $T=13460 52460 0 0 $X=13380 $Y=52050
X32 22 M3_M2_CDNS_765068464212 $T=13460 61710 0 0 $X=13380 $Y=61300
X33 22 M3_M2_CDNS_765068464212 $T=13460 71540 0 0 $X=13380 $Y=71130
X34 1 M3_M2_CDNS_765068464212 $T=33680 34900 0 0 $X=33600 $Y=34490
X35 2 M3_M2_CDNS_765068464212 $T=34530 43540 0 0 $X=34450 $Y=43130
X36 23 M3_M2_CDNS_765068464212 $T=34980 34600 0 0 $X=34900 $Y=34190
X37 19 M3_M2_CDNS_765068464212 $T=35730 51660 0 0 $X=35650 $Y=51250
X38 23 M3_M2_CDNS_765068464212 $T=35830 43240 0 0 $X=35750 $Y=42830
X39 23 M3_M2_CDNS_765068464212 $T=37030 51360 0 0 $X=36950 $Y=50950
X40 20 M3_M2_CDNS_765068464212 $T=37620 59850 0 0 $X=37540 $Y=59440
X41 23 M3_M2_CDNS_765068464212 $T=38920 59550 0 0 $X=38840 $Y=59140
X42 1 M3_M2_CDNS_765068464212 $T=60120 25320 0 0 $X=60040 $Y=24910
X43 2 M3_M2_CDNS_765068464212 $T=60360 34570 0 0 $X=60280 $Y=34160
X44 19 M3_M2_CDNS_765068464212 $T=60910 42670 0 0 $X=60830 $Y=42260
X45 24 M3_M2_CDNS_765068464212 $T=61420 25010 0 0 $X=61340 $Y=24600
X46 24 M3_M2_CDNS_765068464212 $T=61660 34270 0 0 $X=61580 $Y=33860
X47 24 M3_M2_CDNS_765068464212 $T=62210 42370 0 0 $X=62130 $Y=41960
X48 20 M3_M2_CDNS_765068464212 $T=62340 50730 0 0 $X=62260 $Y=50320
X49 24 M3_M2_CDNS_765068464212 $T=63640 50430 0 0 $X=63560 $Y=50020
X50 19 M2_M1_CDNS_765068464213 $T=3540 68870 0 0 $X=3460 $Y=68460
X51 20 M2_M1_CDNS_765068464213 $T=3540 78670 0 0 $X=3460 $Y=78260
X52 1 M2_M1_CDNS_765068464213 $T=3840 48140 0 0 $X=3760 $Y=47730
X53 2 M2_M1_CDNS_765068464213 $T=3840 57600 0 0 $X=3760 $Y=57190
X54 21 M2_M1_CDNS_765068464213 $T=4840 68580 0 0 $X=4760 $Y=68170
X55 21 M2_M1_CDNS_765068464213 $T=4840 78370 0 0 $X=4760 $Y=77960
X56 21 M2_M1_CDNS_765068464213 $T=5140 47840 0 0 $X=5060 $Y=47430
X57 21 M2_M1_CDNS_765068464213 $T=5140 57310 0 0 $X=5060 $Y=56900
X58 1 M2_M1_CDNS_765068464213 $T=12060 42520 0 0 $X=11980 $Y=42110
X59 2 M2_M1_CDNS_765068464213 $T=12160 52760 0 0 $X=12080 $Y=52350
X60 19 M2_M1_CDNS_765068464213 $T=12160 62010 0 0 $X=12080 $Y=61600
X61 20 M2_M1_CDNS_765068464213 $T=12160 71820 0 0 $X=12080 $Y=71410
X62 22 M2_M1_CDNS_765068464213 $T=13360 42210 0 0 $X=13280 $Y=41800
X63 22 M2_M1_CDNS_765068464213 $T=13460 52460 0 0 $X=13380 $Y=52050
X64 22 M2_M1_CDNS_765068464213 $T=13460 61710 0 0 $X=13380 $Y=61300
X65 22 M2_M1_CDNS_765068464213 $T=13460 71540 0 0 $X=13380 $Y=71130
X66 1 M2_M1_CDNS_765068464213 $T=33680 34900 0 0 $X=33600 $Y=34490
X67 2 M2_M1_CDNS_765068464213 $T=34530 43540 0 0 $X=34450 $Y=43130
X68 23 M2_M1_CDNS_765068464213 $T=34980 34600 0 0 $X=34900 $Y=34190
X69 19 M2_M1_CDNS_765068464213 $T=35730 51660 0 0 $X=35650 $Y=51250
X70 23 M2_M1_CDNS_765068464213 $T=35830 43240 0 0 $X=35750 $Y=42830
X71 23 M2_M1_CDNS_765068464213 $T=37030 51360 0 0 $X=36950 $Y=50950
X72 20 M2_M1_CDNS_765068464213 $T=37620 59850 0 0 $X=37540 $Y=59440
X73 23 M2_M1_CDNS_765068464213 $T=38920 59550 0 0 $X=38840 $Y=59140
X74 1 M2_M1_CDNS_765068464213 $T=60120 25320 0 0 $X=60040 $Y=24910
X75 2 M2_M1_CDNS_765068464213 $T=60360 34570 0 0 $X=60280 $Y=34160
X76 19 M2_M1_CDNS_765068464213 $T=60910 42670 0 0 $X=60830 $Y=42260
X77 24 M2_M1_CDNS_765068464213 $T=61420 25010 0 0 $X=61340 $Y=24600
X78 24 M2_M1_CDNS_765068464213 $T=61660 34270 0 0 $X=61580 $Y=33860
X79 24 M2_M1_CDNS_765068464213 $T=62210 42370 0 0 $X=62130 $Y=41960
X80 20 M2_M1_CDNS_765068464213 $T=62340 50730 0 0 $X=62260 $Y=50320
X81 24 M2_M1_CDNS_765068464213 $T=63640 50430 0 0 $X=63560 $Y=50020
X82 19 M4_M3_CDNS_765068464214 $T=550 69610 0 0 $X=110 $Y=69200
X83 20 M4_M3_CDNS_765068464214 $T=740 78860 0 0 $X=300 $Y=78450
X84 25 M4_M3_CDNS_765068464215 $T=8040 45040 0 0 $X=7680 $Y=44910
X85 25 M4_M3_CDNS_765068464215 $T=8040 54400 0 0 $X=7680 $Y=54270
X86 25 M4_M3_CDNS_765068464215 $T=8040 65960 0 0 $X=7680 $Y=65830
X87 25 M4_M3_CDNS_765068464215 $T=8040 75820 0 0 $X=7680 $Y=75690
X88 26 M4_M3_CDNS_765068464215 $T=9700 49570 0 0 $X=9340 $Y=49440
X89 26 M4_M3_CDNS_765068464215 $T=9700 56020 0 0 $X=9340 $Y=55890
X90 26 M4_M3_CDNS_765068464215 $T=9700 70720 0 0 $X=9340 $Y=70590
X91 26 M4_M3_CDNS_765068464215 $T=10210 80980 0 0 $X=9850 $Y=80850
X92 25 M4_M3_CDNS_765068464215 $T=15410 39170 0 0 $X=15050 $Y=39040
X93 25 M4_M3_CDNS_765068464215 $T=15410 49510 0 0 $X=15050 $Y=49380
X94 25 M4_M3_CDNS_765068464215 $T=16420 59350 0 0 $X=16060 $Y=59220
X95 25 M4_M3_CDNS_765068464215 $T=16420 69100 0 0 $X=16060 $Y=68970
X96 26 M4_M3_CDNS_765068464215 $T=20090 46310 0 0 $X=19730 $Y=46180
X97 26 M4_M3_CDNS_765068464215 $T=20090 54850 0 0 $X=19730 $Y=54720
X98 26 M4_M3_CDNS_765068464215 $T=20090 63060 0 0 $X=19730 $Y=62930
X99 26 M4_M3_CDNS_765068464215 $T=20090 73290 0 0 $X=19730 $Y=73160
X100 25 M4_M3_CDNS_765068464215 $T=21880 40430 0 0 $X=21520 $Y=40300
X101 25 M4_M3_CDNS_765068464215 $T=21880 49270 0 0 $X=21520 $Y=49140
X102 25 M4_M3_CDNS_765068464215 $T=21880 56610 0 0 $X=21520 $Y=56480
X103 25 M4_M3_CDNS_765068464215 $T=21880 65140 0 0 $X=21520 $Y=65010
X104 25 M4_M3_CDNS_765068464215 $T=37610 40150 0 0 $X=37250 $Y=40020
X105 25 M4_M3_CDNS_765068464215 $T=37610 47500 0 0 $X=37250 $Y=47370
X106 25 M4_M3_CDNS_765068464215 $T=38430 32280 0 0 $X=38070 $Y=32150
X107 25 M4_M3_CDNS_765068464215 $T=40870 56200 0 0 $X=40510 $Y=56070
X108 26 M4_M3_CDNS_765068464215 $T=42240 37560 0 0 $X=41880 $Y=37430
X109 26 M4_M3_CDNS_765068464215 $T=42240 46080 0 0 $X=41880 $Y=45950
X110 26 M4_M3_CDNS_765068464215 $T=42240 54850 0 0 $X=41880 $Y=54720
X111 26 M4_M3_CDNS_765068464215 $T=42240 63890 0 0 $X=41880 $Y=63760
X112 26 M4_M3_CDNS_765068464215 $T=42240 83140 0 0 $X=41880 $Y=83010
X113 25 M4_M3_CDNS_765068464215 $T=44540 49270 0 0 $X=44180 $Y=49140
X114 25 M4_M3_CDNS_765068464215 $T=47830 32110 0 0 $X=47470 $Y=31980
X115 25 M4_M3_CDNS_765068464215 $T=47830 40320 0 0 $X=47470 $Y=40190
X116 25 M4_M3_CDNS_765068464215 $T=49050 56510 0 0 $X=48690 $Y=56380
X117 25 M4_M3_CDNS_765068464215 $T=64950 31490 0 0 $X=64590 $Y=31360
X118 25 M4_M3_CDNS_765068464215 $T=64950 39420 0 0 $X=64590 $Y=39290
X119 25 M4_M3_CDNS_765068464215 $T=64950 47290 0 0 $X=64590 $Y=47160
X120 25 M4_M3_CDNS_765068464215 $T=65120 23060 0 0 $X=64760 $Y=22930
X121 26 M4_M3_CDNS_765068464215 $T=67370 29860 0 0 $X=67010 $Y=29730
X122 26 M4_M3_CDNS_765068464215 $T=67370 37290 0 0 $X=67010 $Y=37160
X123 26 M4_M3_CDNS_765068464215 $T=67370 46520 0 0 $X=67010 $Y=46390
X124 26 M4_M3_CDNS_765068464215 $T=69160 53660 0 0 $X=68800 $Y=53530
X125 25 M4_M3_CDNS_765068464215 $T=71460 23060 0 0 $X=71100 $Y=22930
X126 25 M4_M3_CDNS_765068464215 $T=71460 31450 0 0 $X=71100 $Y=31320
X127 25 M4_M3_CDNS_765068464215 $T=71460 39840 0 0 $X=71100 $Y=39710
X128 25 M4_M3_CDNS_765068464215 $T=71460 48230 0 0 $X=71100 $Y=48100
X129 27 M4_M3_CDNS_765068464215 $T=91890 5340 0 0 $X=91530 $Y=5210
X130 25 M3_M2_CDNS_765068464216 $T=8040 45040 0 0 $X=7680 $Y=44910
X131 25 M3_M2_CDNS_765068464216 $T=8040 54400 0 0 $X=7680 $Y=54270
X132 25 M3_M2_CDNS_765068464216 $T=8040 65960 0 0 $X=7680 $Y=65830
X133 25 M3_M2_CDNS_765068464216 $T=8040 75820 0 0 $X=7680 $Y=75690
X134 26 M3_M2_CDNS_765068464216 $T=9700 49570 0 0 $X=9340 $Y=49440
X135 26 M3_M2_CDNS_765068464216 $T=9700 56020 0 0 $X=9340 $Y=55890
X136 26 M3_M2_CDNS_765068464216 $T=9700 70720 0 0 $X=9340 $Y=70590
X137 26 M3_M2_CDNS_765068464216 $T=10210 80980 0 0 $X=9850 $Y=80850
X138 25 M3_M2_CDNS_765068464216 $T=15410 39170 0 0 $X=15050 $Y=39040
X139 25 M3_M2_CDNS_765068464216 $T=15410 49510 0 0 $X=15050 $Y=49380
X140 25 M3_M2_CDNS_765068464216 $T=16420 59350 0 0 $X=16060 $Y=59220
X141 25 M3_M2_CDNS_765068464216 $T=16420 69100 0 0 $X=16060 $Y=68970
X142 26 M3_M2_CDNS_765068464216 $T=20090 46310 0 0 $X=19730 $Y=46180
X143 26 M3_M2_CDNS_765068464216 $T=20090 54850 0 0 $X=19730 $Y=54720
X144 26 M3_M2_CDNS_765068464216 $T=20090 63060 0 0 $X=19730 $Y=62930
X145 26 M3_M2_CDNS_765068464216 $T=20090 73290 0 0 $X=19730 $Y=73160
X146 25 M3_M2_CDNS_765068464216 $T=21880 40430 0 0 $X=21520 $Y=40300
X147 25 M3_M2_CDNS_765068464216 $T=21880 49270 0 0 $X=21520 $Y=49140
X148 25 M3_M2_CDNS_765068464216 $T=21880 56610 0 0 $X=21520 $Y=56480
X149 25 M3_M2_CDNS_765068464216 $T=21880 65140 0 0 $X=21520 $Y=65010
X150 25 M3_M2_CDNS_765068464216 $T=37610 40150 0 0 $X=37250 $Y=40020
X151 25 M3_M2_CDNS_765068464216 $T=37610 47500 0 0 $X=37250 $Y=47370
X152 25 M3_M2_CDNS_765068464216 $T=38430 32280 0 0 $X=38070 $Y=32150
X153 25 M3_M2_CDNS_765068464216 $T=40870 56200 0 0 $X=40510 $Y=56070
X154 26 M3_M2_CDNS_765068464216 $T=42240 37560 0 0 $X=41880 $Y=37430
X155 26 M3_M2_CDNS_765068464216 $T=42240 46080 0 0 $X=41880 $Y=45950
X156 26 M3_M2_CDNS_765068464216 $T=42240 54850 0 0 $X=41880 $Y=54720
X157 26 M3_M2_CDNS_765068464216 $T=42240 63890 0 0 $X=41880 $Y=63760
X158 26 M3_M2_CDNS_765068464216 $T=42240 83140 0 0 $X=41880 $Y=83010
X159 25 M3_M2_CDNS_765068464216 $T=44540 49270 0 0 $X=44180 $Y=49140
X160 25 M3_M2_CDNS_765068464216 $T=47830 32110 0 0 $X=47470 $Y=31980
X161 25 M3_M2_CDNS_765068464216 $T=47830 40320 0 0 $X=47470 $Y=40190
X162 25 M3_M2_CDNS_765068464216 $T=49050 56510 0 0 $X=48690 $Y=56380
X163 25 M3_M2_CDNS_765068464216 $T=64950 31490 0 0 $X=64590 $Y=31360
X164 25 M3_M2_CDNS_765068464216 $T=64950 39420 0 0 $X=64590 $Y=39290
X165 25 M3_M2_CDNS_765068464216 $T=64950 47290 0 0 $X=64590 $Y=47160
X166 25 M3_M2_CDNS_765068464216 $T=65120 23060 0 0 $X=64760 $Y=22930
X167 26 M3_M2_CDNS_765068464216 $T=67370 29860 0 0 $X=67010 $Y=29730
X168 26 M3_M2_CDNS_765068464216 $T=67370 37290 0 0 $X=67010 $Y=37160
X169 26 M3_M2_CDNS_765068464216 $T=67370 46520 0 0 $X=67010 $Y=46390
X170 26 M3_M2_CDNS_765068464216 $T=69160 53660 0 0 $X=68800 $Y=53530
X171 25 M3_M2_CDNS_765068464216 $T=71460 23060 0 0 $X=71100 $Y=22930
X172 25 M3_M2_CDNS_765068464216 $T=71460 31450 0 0 $X=71100 $Y=31320
X173 25 M3_M2_CDNS_765068464216 $T=71460 39840 0 0 $X=71100 $Y=39710
X174 25 M3_M2_CDNS_765068464216 $T=71460 48230 0 0 $X=71100 $Y=48100
X175 27 M3_M2_CDNS_765068464216 $T=91890 5340 0 0 $X=91530 $Y=5210
X176 19 M4_M3_CDNS_765068464217 $T=3540 68870 0 0 $X=3460 $Y=68460
X177 20 M4_M3_CDNS_765068464217 $T=3540 78670 0 0 $X=3460 $Y=78260
X178 1 M4_M3_CDNS_765068464217 $T=3840 48140 0 0 $X=3760 $Y=47730
X179 2 M4_M3_CDNS_765068464217 $T=3840 57600 0 0 $X=3760 $Y=57190
X180 1 M4_M3_CDNS_765068464217 $T=12060 42520 0 0 $X=11980 $Y=42110
X181 20 M4_M3_CDNS_765068464217 $T=12150 71810 0 0 $X=12070 $Y=71400
X182 2 M4_M3_CDNS_765068464217 $T=12160 52760 0 0 $X=12080 $Y=52350
X183 19 M4_M3_CDNS_765068464217 $T=12160 62010 0 0 $X=12080 $Y=61600
X184 1 M4_M3_CDNS_765068464217 $T=33680 34900 0 0 $X=33600 $Y=34490
X185 2 M4_M3_CDNS_765068464217 $T=34530 43540 0 0 $X=34450 $Y=43130
X186 19 M4_M3_CDNS_765068464217 $T=35730 51660 0 0 $X=35650 $Y=51250
X187 20 M4_M3_CDNS_765068464217 $T=37620 59850 0 0 $X=37540 $Y=59440
X188 1 M4_M3_CDNS_765068464217 $T=60120 25320 0 0 $X=60040 $Y=24910
X189 2 M4_M3_CDNS_765068464217 $T=60360 34570 0 0 $X=60280 $Y=34160
X190 19 M4_M3_CDNS_765068464217 $T=60910 42670 0 0 $X=60830 $Y=42260
X191 20 M4_M3_CDNS_765068464217 $T=62340 50730 0 0 $X=62260 $Y=50320
X192 1 M5_M4_CDNS_765068464218 $T=33830 48370 0 0 $X=33750 $Y=48240
X193 2 M5_M4_CDNS_765068464218 $T=34690 57170 0 0 $X=34610 $Y=57040
X194 1 M5_M4_CDNS_765068464218 $T=35210 48370 0 0 $X=35130 $Y=48240
X195 19 M5_M4_CDNS_765068464218 $T=36060 69610 0 0 $X=35980 $Y=69480
X196 2 M5_M4_CDNS_765068464218 $T=36620 57170 0 0 $X=36540 $Y=57040
X197 19 M5_M4_CDNS_765068464218 $T=39250 69610 0 0 $X=39170 $Y=69480
X198 28 M5_M4_CDNS_765068464218 $T=59850 67350 0 0 $X=59770 $Y=67220
X199 28 M5_M4_CDNS_765068464218 $T=64530 67360 0 0 $X=64450 $Y=67230
X200 25 M2_M1_CDNS_765068464219 $T=8040 45040 0 0 $X=7680 $Y=44910
X201 25 M2_M1_CDNS_765068464219 $T=8040 54400 0 0 $X=7680 $Y=54270
X202 25 M2_M1_CDNS_765068464219 $T=8040 65960 0 0 $X=7680 $Y=65830
X203 25 M2_M1_CDNS_765068464219 $T=8040 75820 0 0 $X=7680 $Y=75690
X204 26 M2_M1_CDNS_765068464219 $T=9700 49570 0 0 $X=9340 $Y=49440
X205 26 M2_M1_CDNS_765068464219 $T=9700 56020 0 0 $X=9340 $Y=55890
X206 26 M2_M1_CDNS_765068464219 $T=9700 70720 0 0 $X=9340 $Y=70590
X207 26 M2_M1_CDNS_765068464219 $T=10210 80980 0 0 $X=9850 $Y=80850
X208 25 M2_M1_CDNS_765068464219 $T=15410 39170 0 0 $X=15050 $Y=39040
X209 25 M2_M1_CDNS_765068464219 $T=15410 49510 0 0 $X=15050 $Y=49380
X210 25 M2_M1_CDNS_765068464219 $T=16420 59350 0 0 $X=16060 $Y=59220
X211 25 M2_M1_CDNS_765068464219 $T=16420 69100 0 0 $X=16060 $Y=68970
X212 26 M2_M1_CDNS_765068464219 $T=20090 46310 0 0 $X=19730 $Y=46180
X213 26 M2_M1_CDNS_765068464219 $T=20090 54850 0 0 $X=19730 $Y=54720
X214 26 M2_M1_CDNS_765068464219 $T=20090 63060 0 0 $X=19730 $Y=62930
X215 26 M2_M1_CDNS_765068464219 $T=20090 73290 0 0 $X=19730 $Y=73160
X216 25 M2_M1_CDNS_765068464219 $T=21880 40430 0 0 $X=21520 $Y=40300
X217 25 M2_M1_CDNS_765068464219 $T=21880 49270 0 0 $X=21520 $Y=49140
X218 25 M2_M1_CDNS_765068464219 $T=21880 56610 0 0 $X=21520 $Y=56480
X219 25 M2_M1_CDNS_765068464219 $T=21880 65140 0 0 $X=21520 $Y=65010
X220 25 M2_M1_CDNS_765068464219 $T=37610 40150 0 0 $X=37250 $Y=40020
X221 25 M2_M1_CDNS_765068464219 $T=37610 47500 0 0 $X=37250 $Y=47370
X222 25 M2_M1_CDNS_765068464219 $T=38430 32280 0 0 $X=38070 $Y=32150
X223 25 M2_M1_CDNS_765068464219 $T=40870 56200 0 0 $X=40510 $Y=56070
X224 26 M2_M1_CDNS_765068464219 $T=42240 37560 0 0 $X=41880 $Y=37430
X225 26 M2_M1_CDNS_765068464219 $T=42240 46080 0 0 $X=41880 $Y=45950
X226 26 M2_M1_CDNS_765068464219 $T=42240 54850 0 0 $X=41880 $Y=54720
X227 26 M2_M1_CDNS_765068464219 $T=42240 63890 0 0 $X=41880 $Y=63760
X228 26 M2_M1_CDNS_765068464219 $T=42240 83140 0 0 $X=41880 $Y=83010
X229 25 M2_M1_CDNS_765068464219 $T=44540 49270 0 0 $X=44180 $Y=49140
X230 25 M2_M1_CDNS_765068464219 $T=47830 32110 0 0 $X=47470 $Y=31980
X231 25 M2_M1_CDNS_765068464219 $T=47830 40320 0 0 $X=47470 $Y=40190
X232 25 M2_M1_CDNS_765068464219 $T=49050 56510 0 0 $X=48690 $Y=56380
X233 25 M2_M1_CDNS_765068464219 $T=64950 31490 0 0 $X=64590 $Y=31360
X234 25 M2_M1_CDNS_765068464219 $T=64950 39420 0 0 $X=64590 $Y=39290
X235 25 M2_M1_CDNS_765068464219 $T=64950 47290 0 0 $X=64590 $Y=47160
X236 25 M2_M1_CDNS_765068464219 $T=65120 23060 0 0 $X=64760 $Y=22930
X237 26 M2_M1_CDNS_765068464219 $T=67370 29860 0 0 $X=67010 $Y=29730
X238 26 M2_M1_CDNS_765068464219 $T=67370 37290 0 0 $X=67010 $Y=37160
X239 26 M2_M1_CDNS_765068464219 $T=67370 46520 0 0 $X=67010 $Y=46390
X240 26 M2_M1_CDNS_765068464219 $T=69160 53660 0 0 $X=68800 $Y=53530
X241 25 M2_M1_CDNS_765068464219 $T=71460 23060 0 0 $X=71100 $Y=22930
X242 25 M2_M1_CDNS_765068464219 $T=71460 31450 0 0 $X=71100 $Y=31320
X243 25 M2_M1_CDNS_765068464219 $T=71460 39840 0 0 $X=71100 $Y=39710
X244 25 M2_M1_CDNS_765068464219 $T=71460 48230 0 0 $X=71100 $Y=48100
X245 27 M2_M1_CDNS_765068464219 $T=91890 5340 0 0 $X=91530 $Y=5210
X246 29 M4_M3_CDNS_7650684642110 $T=34420 41500 0 0 $X=34340 $Y=41370
X247 30 M4_M3_CDNS_7650684642110 $T=35180 50790 0 0 $X=35100 $Y=50660
X248 31 M4_M3_CDNS_7650684642110 $T=36700 58320 0 0 $X=36620 $Y=58190
X249 28 M4_M3_CDNS_7650684642110 $T=38150 67350 0 0 $X=38070 $Y=67220
X250 29 M4_M3_CDNS_7650684642110 $T=39220 41500 0 0 $X=39140 $Y=41370
X251 30 M4_M3_CDNS_7650684642110 $T=40000 50780 0 0 $X=39920 $Y=50650
X252 31 M4_M3_CDNS_7650684642110 $T=43090 58320 0 0 $X=43010 $Y=58190
X253 32 M4_M3_CDNS_7650684642110 $T=60680 32400 0 0 $X=60600 $Y=32270
X254 33 M4_M3_CDNS_7650684642110 $T=60890 40780 0 0 $X=60810 $Y=40650
X255 34 M4_M3_CDNS_7650684642110 $T=61780 49010 0 0 $X=61700 $Y=48880
X256 35 M4_M3_CDNS_7650684642110 $T=62920 58800 0 0 $X=62840 $Y=58670
X257 32 M4_M3_CDNS_7650684642110 $T=65120 32400 0 0 $X=65040 $Y=32270
X258 33 M4_M3_CDNS_7650684642110 $T=66260 40780 0 0 $X=66180 $Y=40650
X259 34 M4_M3_CDNS_7650684642110 $T=67200 49000 0 0 $X=67120 $Y=48870
X260 35 M4_M3_CDNS_7650684642110 $T=86280 63220 0 0 $X=86200 $Y=63090
X261 28 M4_M3_CDNS_7650684642110 $T=87220 73220 0 0 $X=87140 $Y=73090
X262 7 M3_M2_CDNS_7650684642111 $T=15370 42570 0 0 $X=15290 $Y=42440
X263 36 M3_M2_CDNS_7650684642111 $T=18560 52730 0 0 $X=18480 $Y=52600
X264 37 M3_M2_CDNS_7650684642111 $T=18760 60810 0 0 $X=18680 $Y=60680
X265 10 M3_M2_CDNS_7650684642111 $T=19170 51720 0 0 $X=19090 $Y=51590
X266 5 M3_M2_CDNS_7650684642111 $T=19210 50780 0 0 $X=19130 $Y=50650
X267 6 M3_M2_CDNS_7650684642111 $T=20100 59120 0 0 $X=20020 $Y=58990
X268 8 M3_M2_CDNS_7650684642111 $T=20110 60060 0 0 $X=20030 $Y=59930
X269 38 M3_M2_CDNS_7650684642111 $T=21310 44360 0 0 $X=21230 $Y=44230
X270 9 M3_M2_CDNS_7650684642111 $T=22540 68220 0 0 $X=22460 $Y=68090
X271 3 M3_M2_CDNS_7650684642111 $T=22550 67750 0 0 $X=22470 $Y=67620
X272 12 M3_M2_CDNS_7650684642111 $T=39390 43590 0 0 $X=39310 $Y=43460
X273 11 M3_M2_CDNS_7650684642111 $T=39400 34950 0 0 $X=39320 $Y=34820
X274 39 M3_M2_CDNS_7650684642111 $T=40580 34370 0 0 $X=40500 $Y=34240
X275 13 M3_M2_CDNS_7650684642111 $T=41300 51720 0 0 $X=41220 $Y=51590
X276 14 M3_M2_CDNS_7650684642111 $T=43140 59910 0 0 $X=43060 $Y=59780
X277 40 M3_M2_CDNS_7650684642111 $T=44180 43130 0 0 $X=44100 $Y=43000
X278 41 M3_M2_CDNS_7650684642111 $T=44260 51280 0 0 $X=44180 $Y=51150
X279 42 M3_M2_CDNS_7650684642111 $T=44310 34880 0 0 $X=44230 $Y=34750
X280 16 M3_M2_CDNS_7650684642111 $T=66170 34680 0 0 $X=66090 $Y=34550
X281 15 M3_M2_CDNS_7650684642111 $T=66360 26140 0 0 $X=66280 $Y=26010
X282 17 M3_M2_CDNS_7650684642111 $T=66510 43080 0 0 $X=66430 $Y=42950
X283 43 M3_M2_CDNS_7650684642111 $T=67390 25350 0 0 $X=67310 $Y=25220
X284 18 M3_M2_CDNS_7650684642111 $T=68160 51630 0 0 $X=68080 $Y=51500
X285 44 M3_M2_CDNS_7650684642111 $T=69560 42730 0 0 $X=69480 $Y=42600
X286 45 M3_M2_CDNS_7650684642111 $T=69650 25880 0 0 $X=69570 $Y=25750
X287 46 M3_M2_CDNS_7650684642111 $T=69930 34320 0 0 $X=69850 $Y=34190
X288 25 M5_M4_CDNS_7650684642113 $T=8040 45040 0 0 $X=7680 $Y=44910
X289 25 M5_M4_CDNS_7650684642113 $T=8040 54400 0 0 $X=7680 $Y=54270
X290 25 M5_M4_CDNS_7650684642113 $T=8040 65960 0 0 $X=7680 $Y=65830
X291 25 M5_M4_CDNS_7650684642113 $T=8040 75820 0 0 $X=7680 $Y=75690
X292 26 M5_M4_CDNS_7650684642113 $T=9700 49570 0 0 $X=9340 $Y=49440
X293 26 M5_M4_CDNS_7650684642113 $T=9700 56020 0 0 $X=9340 $Y=55890
X294 26 M5_M4_CDNS_7650684642113 $T=9700 70720 0 0 $X=9340 $Y=70590
X295 26 M5_M4_CDNS_7650684642113 $T=10210 80980 0 0 $X=9850 $Y=80850
X296 25 M5_M4_CDNS_7650684642113 $T=15410 39170 0 0 $X=15050 $Y=39040
X297 25 M5_M4_CDNS_7650684642113 $T=15410 49510 0 0 $X=15050 $Y=49380
X298 25 M5_M4_CDNS_7650684642113 $T=16420 59350 0 0 $X=16060 $Y=59220
X299 25 M5_M4_CDNS_7650684642113 $T=16420 69100 0 0 $X=16060 $Y=68970
X300 26 M5_M4_CDNS_7650684642113 $T=20090 46310 0 0 $X=19730 $Y=46180
X301 26 M5_M4_CDNS_7650684642113 $T=20090 54850 0 0 $X=19730 $Y=54720
X302 26 M5_M4_CDNS_7650684642113 $T=20090 63060 0 0 $X=19730 $Y=62930
X303 26 M5_M4_CDNS_7650684642113 $T=20090 73290 0 0 $X=19730 $Y=73160
X304 25 M5_M4_CDNS_7650684642113 $T=21880 40430 0 0 $X=21520 $Y=40300
X305 25 M5_M4_CDNS_7650684642113 $T=21880 49270 0 0 $X=21520 $Y=49140
X306 25 M5_M4_CDNS_7650684642113 $T=21880 56610 0 0 $X=21520 $Y=56480
X307 25 M5_M4_CDNS_7650684642113 $T=21880 65140 0 0 $X=21520 $Y=65010
X308 25 M5_M4_CDNS_7650684642113 $T=37610 40150 0 0 $X=37250 $Y=40020
X309 25 M5_M4_CDNS_7650684642113 $T=37610 47500 0 0 $X=37250 $Y=47370
X310 25 M5_M4_CDNS_7650684642113 $T=38430 32280 0 0 $X=38070 $Y=32150
X311 25 M5_M4_CDNS_7650684642113 $T=40870 56200 0 0 $X=40510 $Y=56070
X312 26 M5_M4_CDNS_7650684642113 $T=42240 37560 0 0 $X=41880 $Y=37430
X313 26 M5_M4_CDNS_7650684642113 $T=42240 46080 0 0 $X=41880 $Y=45950
X314 26 M5_M4_CDNS_7650684642113 $T=42240 54850 0 0 $X=41880 $Y=54720
X315 26 M5_M4_CDNS_7650684642113 $T=42240 63890 0 0 $X=41880 $Y=63760
X316 26 M5_M4_CDNS_7650684642113 $T=42240 83140 0 0 $X=41880 $Y=83010
X317 25 M5_M4_CDNS_7650684642113 $T=44540 49270 0 0 $X=44180 $Y=49140
X318 25 M5_M4_CDNS_7650684642113 $T=47830 32110 0 0 $X=47470 $Y=31980
X319 25 M5_M4_CDNS_7650684642113 $T=47830 40320 0 0 $X=47470 $Y=40190
X320 25 M5_M4_CDNS_7650684642113 $T=49050 56510 0 0 $X=48690 $Y=56380
X321 25 M5_M4_CDNS_7650684642113 $T=64950 31490 0 0 $X=64590 $Y=31360
X322 25 M5_M4_CDNS_7650684642113 $T=64950 39420 0 0 $X=64590 $Y=39290
X323 25 M5_M4_CDNS_7650684642113 $T=64950 47290 0 0 $X=64590 $Y=47160
X324 25 M5_M4_CDNS_7650684642113 $T=65120 23060 0 0 $X=64760 $Y=22930
X325 26 M5_M4_CDNS_7650684642113 $T=67370 29860 0 0 $X=67010 $Y=29730
X326 26 M5_M4_CDNS_7650684642113 $T=67370 37290 0 0 $X=67010 $Y=37160
X327 26 M5_M4_CDNS_7650684642113 $T=67370 46520 0 0 $X=67010 $Y=46390
X328 26 M5_M4_CDNS_7650684642113 $T=69160 53660 0 0 $X=68800 $Y=53530
X329 25 M5_M4_CDNS_7650684642113 $T=71460 23060 0 0 $X=71100 $Y=22930
X330 25 M5_M4_CDNS_7650684642113 $T=71460 31450 0 0 $X=71100 $Y=31320
X331 25 M5_M4_CDNS_7650684642113 $T=71460 39840 0 0 $X=71100 $Y=39710
X332 25 M5_M4_CDNS_7650684642113 $T=71460 48230 0 0 $X=71100 $Y=48100
X333 27 M5_M4_CDNS_7650684642113 $T=91890 5340 0 0 $X=91530 $Y=5210
X334 25 M6_M5_CDNS_7650684642114 $T=8040 45040 0 0 $X=7680 $Y=44910
X335 25 M6_M5_CDNS_7650684642114 $T=8040 54400 0 0 $X=7680 $Y=54270
X336 25 M6_M5_CDNS_7650684642114 $T=8040 65960 0 0 $X=7680 $Y=65830
X337 25 M6_M5_CDNS_7650684642114 $T=8040 75820 0 0 $X=7680 $Y=75690
X338 26 M6_M5_CDNS_7650684642114 $T=9700 49570 0 0 $X=9340 $Y=49440
X339 26 M6_M5_CDNS_7650684642114 $T=9700 56020 0 0 $X=9340 $Y=55890
X340 26 M6_M5_CDNS_7650684642114 $T=9700 70720 0 0 $X=9340 $Y=70590
X341 26 M6_M5_CDNS_7650684642114 $T=10210 80980 0 0 $X=9850 $Y=80850
X342 25 M6_M5_CDNS_7650684642114 $T=15410 39170 0 0 $X=15050 $Y=39040
X343 25 M6_M5_CDNS_7650684642114 $T=15410 49510 0 0 $X=15050 $Y=49380
X344 25 M6_M5_CDNS_7650684642114 $T=16420 59350 0 0 $X=16060 $Y=59220
X345 25 M6_M5_CDNS_7650684642114 $T=16420 69100 0 0 $X=16060 $Y=68970
X346 26 M6_M5_CDNS_7650684642114 $T=20090 46310 0 0 $X=19730 $Y=46180
X347 26 M6_M5_CDNS_7650684642114 $T=20090 54850 0 0 $X=19730 $Y=54720
X348 26 M6_M5_CDNS_7650684642114 $T=20090 63060 0 0 $X=19730 $Y=62930
X349 26 M6_M5_CDNS_7650684642114 $T=20090 73290 0 0 $X=19730 $Y=73160
X350 25 M6_M5_CDNS_7650684642114 $T=21880 40430 0 0 $X=21520 $Y=40300
X351 25 M6_M5_CDNS_7650684642114 $T=21880 49270 0 0 $X=21520 $Y=49140
X352 25 M6_M5_CDNS_7650684642114 $T=21880 56610 0 0 $X=21520 $Y=56480
X353 25 M6_M5_CDNS_7650684642114 $T=21880 65140 0 0 $X=21520 $Y=65010
X354 25 M6_M5_CDNS_7650684642114 $T=37610 40150 0 0 $X=37250 $Y=40020
X355 25 M6_M5_CDNS_7650684642114 $T=37610 47500 0 0 $X=37250 $Y=47370
X356 25 M6_M5_CDNS_7650684642114 $T=38430 32280 0 0 $X=38070 $Y=32150
X357 25 M6_M5_CDNS_7650684642114 $T=40870 56200 0 0 $X=40510 $Y=56070
X358 26 M6_M5_CDNS_7650684642114 $T=42240 37560 0 0 $X=41880 $Y=37430
X359 26 M6_M5_CDNS_7650684642114 $T=42240 46080 0 0 $X=41880 $Y=45950
X360 26 M6_M5_CDNS_7650684642114 $T=42240 54850 0 0 $X=41880 $Y=54720
X361 26 M6_M5_CDNS_7650684642114 $T=42240 63890 0 0 $X=41880 $Y=63760
X362 26 M6_M5_CDNS_7650684642114 $T=42240 83140 0 0 $X=41880 $Y=83010
X363 25 M6_M5_CDNS_7650684642114 $T=44540 49270 0 0 $X=44180 $Y=49140
X364 25 M6_M5_CDNS_7650684642114 $T=47830 32110 0 0 $X=47470 $Y=31980
X365 25 M6_M5_CDNS_7650684642114 $T=47830 40320 0 0 $X=47470 $Y=40190
X366 25 M6_M5_CDNS_7650684642114 $T=49050 56510 0 0 $X=48690 $Y=56380
X367 25 M6_M5_CDNS_7650684642114 $T=64950 31490 0 0 $X=64590 $Y=31360
X368 25 M6_M5_CDNS_7650684642114 $T=64950 39420 0 0 $X=64590 $Y=39290
X369 25 M6_M5_CDNS_7650684642114 $T=64950 47290 0 0 $X=64590 $Y=47160
X370 25 M6_M5_CDNS_7650684642114 $T=65120 23060 0 0 $X=64760 $Y=22930
X371 26 M6_M5_CDNS_7650684642114 $T=67370 29860 0 0 $X=67010 $Y=29730
X372 26 M6_M5_CDNS_7650684642114 $T=67370 37290 0 0 $X=67010 $Y=37160
X373 26 M6_M5_CDNS_7650684642114 $T=67370 46520 0 0 $X=67010 $Y=46390
X374 26 M6_M5_CDNS_7650684642114 $T=69160 53660 0 0 $X=68800 $Y=53530
X375 25 M6_M5_CDNS_7650684642114 $T=71460 23060 0 0 $X=71100 $Y=22930
X376 25 M6_M5_CDNS_7650684642114 $T=71460 31450 0 0 $X=71100 $Y=31320
X377 25 M6_M5_CDNS_7650684642114 $T=71460 39840 0 0 $X=71100 $Y=39710
X378 25 M6_M5_CDNS_7650684642114 $T=71460 48230 0 0 $X=71100 $Y=48100
X379 27 M6_M5_CDNS_7650684642114 $T=91890 5340 0 0 $X=91530 $Y=5210
X380 25 M7_M6_CDNS_7650684642115 $T=8040 45040 0 0 $X=7680 $Y=44910
X381 25 M7_M6_CDNS_7650684642115 $T=8040 54400 0 0 $X=7680 $Y=54270
X382 25 M7_M6_CDNS_7650684642115 $T=8040 65960 0 0 $X=7680 $Y=65830
X383 25 M7_M6_CDNS_7650684642115 $T=8040 75820 0 0 $X=7680 $Y=75690
X384 26 M7_M6_CDNS_7650684642115 $T=9700 49570 0 0 $X=9340 $Y=49440
X385 26 M7_M6_CDNS_7650684642115 $T=9700 56020 0 0 $X=9340 $Y=55890
X386 26 M7_M6_CDNS_7650684642115 $T=9700 70720 0 0 $X=9340 $Y=70590
X387 26 M7_M6_CDNS_7650684642115 $T=10210 80980 0 0 $X=9850 $Y=80850
X388 25 M7_M6_CDNS_7650684642115 $T=15410 39170 0 0 $X=15050 $Y=39040
X389 25 M7_M6_CDNS_7650684642115 $T=15410 49510 0 0 $X=15050 $Y=49380
X390 25 M7_M6_CDNS_7650684642115 $T=16420 59350 0 0 $X=16060 $Y=59220
X391 25 M7_M6_CDNS_7650684642115 $T=16420 69100 0 0 $X=16060 $Y=68970
X392 26 M7_M6_CDNS_7650684642115 $T=20090 46310 0 0 $X=19730 $Y=46180
X393 26 M7_M6_CDNS_7650684642115 $T=20090 54850 0 0 $X=19730 $Y=54720
X394 26 M7_M6_CDNS_7650684642115 $T=20090 63060 0 0 $X=19730 $Y=62930
X395 26 M7_M6_CDNS_7650684642115 $T=20090 73290 0 0 $X=19730 $Y=73160
X396 25 M7_M6_CDNS_7650684642115 $T=21880 40430 0 0 $X=21520 $Y=40300
X397 25 M7_M6_CDNS_7650684642115 $T=21880 49270 0 0 $X=21520 $Y=49140
X398 25 M7_M6_CDNS_7650684642115 $T=21880 56610 0 0 $X=21520 $Y=56480
X399 25 M7_M6_CDNS_7650684642115 $T=21880 65140 0 0 $X=21520 $Y=65010
X400 25 M7_M6_CDNS_7650684642115 $T=37610 40150 0 0 $X=37250 $Y=40020
X401 25 M7_M6_CDNS_7650684642115 $T=37610 47500 0 0 $X=37250 $Y=47370
X402 25 M7_M6_CDNS_7650684642115 $T=38430 32280 0 0 $X=38070 $Y=32150
X403 25 M7_M6_CDNS_7650684642115 $T=40870 56200 0 0 $X=40510 $Y=56070
X404 26 M7_M6_CDNS_7650684642115 $T=42240 37560 0 0 $X=41880 $Y=37430
X405 26 M7_M6_CDNS_7650684642115 $T=42240 46080 0 0 $X=41880 $Y=45950
X406 26 M7_M6_CDNS_7650684642115 $T=42240 54850 0 0 $X=41880 $Y=54720
X407 26 M7_M6_CDNS_7650684642115 $T=42240 63890 0 0 $X=41880 $Y=63760
X408 26 M7_M6_CDNS_7650684642115 $T=42240 83140 0 0 $X=41880 $Y=83010
X409 25 M7_M6_CDNS_7650684642115 $T=44540 49270 0 0 $X=44180 $Y=49140
X410 25 M7_M6_CDNS_7650684642115 $T=47830 32110 0 0 $X=47470 $Y=31980
X411 25 M7_M6_CDNS_7650684642115 $T=47830 40320 0 0 $X=47470 $Y=40190
X412 25 M7_M6_CDNS_7650684642115 $T=49050 56510 0 0 $X=48690 $Y=56380
X413 25 M7_M6_CDNS_7650684642115 $T=64950 31490 0 0 $X=64590 $Y=31360
X414 25 M7_M6_CDNS_7650684642115 $T=64950 39420 0 0 $X=64590 $Y=39290
X415 25 M7_M6_CDNS_7650684642115 $T=64950 47290 0 0 $X=64590 $Y=47160
X416 25 M7_M6_CDNS_7650684642115 $T=65120 23060 0 0 $X=64760 $Y=22930
X417 26 M7_M6_CDNS_7650684642115 $T=67370 29860 0 0 $X=67010 $Y=29730
X418 26 M7_M6_CDNS_7650684642115 $T=67370 37290 0 0 $X=67010 $Y=37160
X419 26 M7_M6_CDNS_7650684642115 $T=67370 46520 0 0 $X=67010 $Y=46390
X420 26 M7_M6_CDNS_7650684642115 $T=69160 53660 0 0 $X=68800 $Y=53530
X421 25 M7_M6_CDNS_7650684642115 $T=71460 23060 0 0 $X=71100 $Y=22930
X422 25 M7_M6_CDNS_7650684642115 $T=71460 31450 0 0 $X=71100 $Y=31320
X423 25 M7_M6_CDNS_7650684642115 $T=71460 39840 0 0 $X=71100 $Y=39710
X424 25 M7_M6_CDNS_7650684642115 $T=71460 48230 0 0 $X=71100 $Y=48100
X425 27 M7_M6_CDNS_7650684642115 $T=91890 5340 0 0 $X=91530 $Y=5210
X426 25 M8_M7_CDNS_7650684642116 $T=8040 45040 0 0 $X=7680 $Y=44910
X427 25 M8_M7_CDNS_7650684642116 $T=8040 54400 0 0 $X=7680 $Y=54270
X428 25 M8_M7_CDNS_7650684642116 $T=8040 65960 0 0 $X=7680 $Y=65830
X429 25 M8_M7_CDNS_7650684642116 $T=8040 75820 0 0 $X=7680 $Y=75690
X430 26 M8_M7_CDNS_7650684642116 $T=9700 49570 0 0 $X=9340 $Y=49440
X431 26 M8_M7_CDNS_7650684642116 $T=9700 56020 0 0 $X=9340 $Y=55890
X432 26 M8_M7_CDNS_7650684642116 $T=9700 70720 0 0 $X=9340 $Y=70590
X433 26 M8_M7_CDNS_7650684642116 $T=10210 80980 0 0 $X=9850 $Y=80850
X434 25 M8_M7_CDNS_7650684642116 $T=15410 39170 0 0 $X=15050 $Y=39040
X435 25 M8_M7_CDNS_7650684642116 $T=15410 49510 0 0 $X=15050 $Y=49380
X436 25 M8_M7_CDNS_7650684642116 $T=16420 59350 0 0 $X=16060 $Y=59220
X437 25 M8_M7_CDNS_7650684642116 $T=16420 69100 0 0 $X=16060 $Y=68970
X438 26 M8_M7_CDNS_7650684642116 $T=20090 46310 0 0 $X=19730 $Y=46180
X439 26 M8_M7_CDNS_7650684642116 $T=20090 54850 0 0 $X=19730 $Y=54720
X440 26 M8_M7_CDNS_7650684642116 $T=20090 63060 0 0 $X=19730 $Y=62930
X441 26 M8_M7_CDNS_7650684642116 $T=20090 73290 0 0 $X=19730 $Y=73160
X442 25 M8_M7_CDNS_7650684642116 $T=21880 40430 0 0 $X=21520 $Y=40300
X443 25 M8_M7_CDNS_7650684642116 $T=21880 49270 0 0 $X=21520 $Y=49140
X444 25 M8_M7_CDNS_7650684642116 $T=21880 56610 0 0 $X=21520 $Y=56480
X445 25 M8_M7_CDNS_7650684642116 $T=21880 65140 0 0 $X=21520 $Y=65010
X446 25 M8_M7_CDNS_7650684642116 $T=37610 40150 0 0 $X=37250 $Y=40020
X447 25 M8_M7_CDNS_7650684642116 $T=37610 47500 0 0 $X=37250 $Y=47370
X448 25 M8_M7_CDNS_7650684642116 $T=38430 32280 0 0 $X=38070 $Y=32150
X449 25 M8_M7_CDNS_7650684642116 $T=40870 56200 0 0 $X=40510 $Y=56070
X450 26 M8_M7_CDNS_7650684642116 $T=42240 37560 0 0 $X=41880 $Y=37430
X451 26 M8_M7_CDNS_7650684642116 $T=42240 46080 0 0 $X=41880 $Y=45950
X452 26 M8_M7_CDNS_7650684642116 $T=42240 54850 0 0 $X=41880 $Y=54720
X453 26 M8_M7_CDNS_7650684642116 $T=42240 63890 0 0 $X=41880 $Y=63760
X454 26 M8_M7_CDNS_7650684642116 $T=42240 83140 0 0 $X=41880 $Y=83010
X455 25 M8_M7_CDNS_7650684642116 $T=44540 49270 0 0 $X=44180 $Y=49140
X456 25 M8_M7_CDNS_7650684642116 $T=47830 32110 0 0 $X=47470 $Y=31980
X457 25 M8_M7_CDNS_7650684642116 $T=47830 40320 0 0 $X=47470 $Y=40190
X458 25 M8_M7_CDNS_7650684642116 $T=49050 56510 0 0 $X=48690 $Y=56380
X459 25 M8_M7_CDNS_7650684642116 $T=64950 31490 0 0 $X=64590 $Y=31360
X460 25 M8_M7_CDNS_7650684642116 $T=64950 39420 0 0 $X=64590 $Y=39290
X461 25 M8_M7_CDNS_7650684642116 $T=64950 47290 0 0 $X=64590 $Y=47160
X462 25 M8_M7_CDNS_7650684642116 $T=65120 23060 0 0 $X=64760 $Y=22930
X463 26 M8_M7_CDNS_7650684642116 $T=67370 29860 0 0 $X=67010 $Y=29730
X464 26 M8_M7_CDNS_7650684642116 $T=67370 37290 0 0 $X=67010 $Y=37160
X465 26 M8_M7_CDNS_7650684642116 $T=67370 46520 0 0 $X=67010 $Y=46390
X466 26 M8_M7_CDNS_7650684642116 $T=69160 53660 0 0 $X=68800 $Y=53530
X467 25 M8_M7_CDNS_7650684642116 $T=71460 23060 0 0 $X=71100 $Y=22930
X468 25 M8_M7_CDNS_7650684642116 $T=71460 31450 0 0 $X=71100 $Y=31320
X469 25 M8_M7_CDNS_7650684642116 $T=71460 39840 0 0 $X=71100 $Y=39710
X470 25 M8_M7_CDNS_7650684642116 $T=71460 48230 0 0 $X=71100 $Y=48100
X471 27 M8_M7_CDNS_7650684642116 $T=91890 5340 0 0 $X=91530 $Y=5210
X472 25 M9_M8_CDNS_7650684642117 $T=8040 45040 0 0 $X=7680 $Y=44910
X473 25 M9_M8_CDNS_7650684642117 $T=8040 54400 0 0 $X=7680 $Y=54270
X474 25 M9_M8_CDNS_7650684642117 $T=8040 65960 0 0 $X=7680 $Y=65830
X475 25 M9_M8_CDNS_7650684642117 $T=8040 75820 0 0 $X=7680 $Y=75690
X476 26 M9_M8_CDNS_7650684642117 $T=9700 49570 0 0 $X=9340 $Y=49440
X477 26 M9_M8_CDNS_7650684642117 $T=9700 56020 0 0 $X=9340 $Y=55890
X478 26 M9_M8_CDNS_7650684642117 $T=9700 70720 0 0 $X=9340 $Y=70590
X479 26 M9_M8_CDNS_7650684642117 $T=10210 80980 0 0 $X=9850 $Y=80850
X480 25 M9_M8_CDNS_7650684642117 $T=15410 39170 0 0 $X=15050 $Y=39040
X481 25 M9_M8_CDNS_7650684642117 $T=15410 49510 0 0 $X=15050 $Y=49380
X482 25 M9_M8_CDNS_7650684642117 $T=16420 59350 0 0 $X=16060 $Y=59220
X483 25 M9_M8_CDNS_7650684642117 $T=16420 69100 0 0 $X=16060 $Y=68970
X484 26 M9_M8_CDNS_7650684642117 $T=20090 46310 0 0 $X=19730 $Y=46180
X485 26 M9_M8_CDNS_7650684642117 $T=20090 54850 0 0 $X=19730 $Y=54720
X486 26 M9_M8_CDNS_7650684642117 $T=20090 63060 0 0 $X=19730 $Y=62930
X487 26 M9_M8_CDNS_7650684642117 $T=20090 73290 0 0 $X=19730 $Y=73160
X488 25 M9_M8_CDNS_7650684642117 $T=21880 40430 0 0 $X=21520 $Y=40300
X489 25 M9_M8_CDNS_7650684642117 $T=21880 49270 0 0 $X=21520 $Y=49140
X490 25 M9_M8_CDNS_7650684642117 $T=21880 56610 0 0 $X=21520 $Y=56480
X491 25 M9_M8_CDNS_7650684642117 $T=21880 65140 0 0 $X=21520 $Y=65010
X492 25 M9_M8_CDNS_7650684642117 $T=37610 40150 0 0 $X=37250 $Y=40020
X493 25 M9_M8_CDNS_7650684642117 $T=37610 47500 0 0 $X=37250 $Y=47370
X494 25 M9_M8_CDNS_7650684642117 $T=38430 32280 0 0 $X=38070 $Y=32150
X495 25 M9_M8_CDNS_7650684642117 $T=40870 56200 0 0 $X=40510 $Y=56070
X496 26 M9_M8_CDNS_7650684642117 $T=42240 37560 0 0 $X=41880 $Y=37430
X497 26 M9_M8_CDNS_7650684642117 $T=42240 46080 0 0 $X=41880 $Y=45950
X498 26 M9_M8_CDNS_7650684642117 $T=42240 54850 0 0 $X=41880 $Y=54720
X499 26 M9_M8_CDNS_7650684642117 $T=42240 63890 0 0 $X=41880 $Y=63760
X500 26 M9_M8_CDNS_7650684642117 $T=42240 83140 0 0 $X=41880 $Y=83010
X501 25 M9_M8_CDNS_7650684642117 $T=44540 49270 0 0 $X=44180 $Y=49140
X502 25 M9_M8_CDNS_7650684642117 $T=47830 32110 0 0 $X=47470 $Y=31980
X503 25 M9_M8_CDNS_7650684642117 $T=47830 40320 0 0 $X=47470 $Y=40190
X504 25 M9_M8_CDNS_7650684642117 $T=49050 56510 0 0 $X=48690 $Y=56380
X505 25 M9_M8_CDNS_7650684642117 $T=64950 31490 0 0 $X=64590 $Y=31360
X506 25 M9_M8_CDNS_7650684642117 $T=64950 39420 0 0 $X=64590 $Y=39290
X507 25 M9_M8_CDNS_7650684642117 $T=64950 47290 0 0 $X=64590 $Y=47160
X508 25 M9_M8_CDNS_7650684642117 $T=65120 23060 0 0 $X=64760 $Y=22930
X509 26 M9_M8_CDNS_7650684642117 $T=67370 29860 0 0 $X=67010 $Y=29730
X510 26 M9_M8_CDNS_7650684642117 $T=67370 37290 0 0 $X=67010 $Y=37160
X511 26 M9_M8_CDNS_7650684642117 $T=67370 46520 0 0 $X=67010 $Y=46390
X512 26 M9_M8_CDNS_7650684642117 $T=69160 53660 0 0 $X=68800 $Y=53530
X513 25 M9_M8_CDNS_7650684642117 $T=71460 23060 0 0 $X=71100 $Y=22930
X514 25 M9_M8_CDNS_7650684642117 $T=71460 31450 0 0 $X=71100 $Y=31320
X515 25 M9_M8_CDNS_7650684642117 $T=71460 39840 0 0 $X=71100 $Y=39710
X516 25 M9_M8_CDNS_7650684642117 $T=71460 48230 0 0 $X=71100 $Y=48100
X517 27 M9_M8_CDNS_7650684642117 $T=91890 5340 0 0 $X=91530 $Y=5210
X518 25 M10_M9_CDNS_7650684642118 $T=8040 45030 0 0 $X=7080 $Y=44750
X519 25 M10_M9_CDNS_7650684642118 $T=8040 54390 0 0 $X=7080 $Y=54110
X520 25 M10_M9_CDNS_7650684642118 $T=8040 65950 0 0 $X=7080 $Y=65670
X521 25 M10_M9_CDNS_7650684642118 $T=8040 75810 0 0 $X=7080 $Y=75530
X522 26 M10_M9_CDNS_7650684642118 $T=9700 49570 0 0 $X=8740 $Y=49290
X523 26 M10_M9_CDNS_7650684642118 $T=9700 56020 0 0 $X=8740 $Y=55740
X524 26 M10_M9_CDNS_7650684642118 $T=9700 70720 0 0 $X=8740 $Y=70440
X525 26 M10_M9_CDNS_7650684642118 $T=10210 80980 0 0 $X=9250 $Y=80700
X526 25 M10_M9_CDNS_7650684642118 $T=15410 39160 0 0 $X=14450 $Y=38880
X527 25 M10_M9_CDNS_7650684642118 $T=15410 49500 0 0 $X=14450 $Y=49220
X528 25 M10_M9_CDNS_7650684642118 $T=16420 59340 0 0 $X=15460 $Y=59060
X529 25 M10_M9_CDNS_7650684642118 $T=16420 69090 0 0 $X=15460 $Y=68810
X530 26 M10_M9_CDNS_7650684642118 $T=20090 46310 0 0 $X=19130 $Y=46030
X531 26 M10_M9_CDNS_7650684642118 $T=20090 54850 0 0 $X=19130 $Y=54570
X532 26 M10_M9_CDNS_7650684642118 $T=20090 63060 0 0 $X=19130 $Y=62780
X533 26 M10_M9_CDNS_7650684642118 $T=20090 73290 0 0 $X=19130 $Y=73010
X534 25 M10_M9_CDNS_7650684642118 $T=21880 40420 0 0 $X=20920 $Y=40140
X535 25 M10_M9_CDNS_7650684642118 $T=21880 49260 0 0 $X=20920 $Y=48980
X536 25 M10_M9_CDNS_7650684642118 $T=21880 56600 0 0 $X=20920 $Y=56320
X537 25 M10_M9_CDNS_7650684642118 $T=21880 65130 0 0 $X=20920 $Y=64850
X538 25 M10_M9_CDNS_7650684642118 $T=37610 40140 0 0 $X=36650 $Y=39860
X539 25 M10_M9_CDNS_7650684642118 $T=37610 47490 0 0 $X=36650 $Y=47210
X540 25 M10_M9_CDNS_7650684642118 $T=38430 32280 0 0 $X=37470 $Y=32000
X541 25 M10_M9_CDNS_7650684642118 $T=40560 14790 0 0 $X=39600 $Y=14510
X542 25 M10_M9_CDNS_7650684642118 $T=40800 56230 0 0 $X=39840 $Y=55950
X543 26 M10_M9_CDNS_7650684642118 $T=42240 37560 0 0 $X=41280 $Y=37280
X544 26 M10_M9_CDNS_7650684642118 $T=42240 46080 0 0 $X=41280 $Y=45800
X545 26 M10_M9_CDNS_7650684642118 $T=42240 54850 0 0 $X=41280 $Y=54570
X546 26 M10_M9_CDNS_7650684642118 $T=42240 63890 0 0 $X=41280 $Y=63610
X547 26 M10_M9_CDNS_7650684642118 $T=42240 83140 0 0 $X=41280 $Y=82860
X548 25 M10_M9_CDNS_7650684642118 $T=44550 49280 0 0 $X=43590 $Y=49000
X549 25 M10_M9_CDNS_7650684642118 $T=47830 32150 0 0 $X=46870 $Y=31870
X550 25 M10_M9_CDNS_7650684642118 $T=47830 40360 0 0 $X=46870 $Y=40080
X551 25 M10_M9_CDNS_7650684642118 $T=49050 56500 0 0 $X=48090 $Y=56220
X552 25 M10_M9_CDNS_7650684642118 $T=64950 31530 0 0 $X=63990 $Y=31250
X553 25 M10_M9_CDNS_7650684642118 $T=64950 39460 0 0 $X=63990 $Y=39180
X554 25 M10_M9_CDNS_7650684642118 $T=64950 47330 0 0 $X=63990 $Y=47050
X555 25 M10_M9_CDNS_7650684642118 $T=65120 23100 0 0 $X=64160 $Y=22820
X556 26 M10_M9_CDNS_7650684642118 $T=67370 29860 0 0 $X=66410 $Y=29580
X557 26 M10_M9_CDNS_7650684642118 $T=67370 37290 0 0 $X=66410 $Y=37010
X558 26 M10_M9_CDNS_7650684642118 $T=67370 46520 0 0 $X=66410 $Y=46240
X559 26 M10_M9_CDNS_7650684642118 $T=69160 53660 0 0 $X=68200 $Y=53380
X560 25 M10_M9_CDNS_7650684642118 $T=71460 23100 0 0 $X=70500 $Y=22820
X561 25 M10_M9_CDNS_7650684642118 $T=71460 31490 0 0 $X=70500 $Y=31210
X562 25 M10_M9_CDNS_7650684642118 $T=71460 39880 0 0 $X=70500 $Y=39600
X563 25 M10_M9_CDNS_7650684642118 $T=71460 48270 0 0 $X=70500 $Y=47990
X564 27 M10_M9_CDNS_7650684642118 $T=91890 5340 0 0 $X=90930 $Y=5060
X565 26 M11_M10_CDNS_7650684642119 $T=9700 49570 0 0 $X=8740 $Y=49290
X566 26 M11_M10_CDNS_7650684642119 $T=9700 56020 0 0 $X=8740 $Y=55740
X567 26 M11_M10_CDNS_7650684642119 $T=9700 70720 0 0 $X=8740 $Y=70440
X568 26 M11_M10_CDNS_7650684642119 $T=10210 80980 0 0 $X=9250 $Y=80700
X569 26 M11_M10_CDNS_7650684642119 $T=20090 46310 0 0 $X=19130 $Y=46030
X570 26 M11_M10_CDNS_7650684642119 $T=20090 54850 0 0 $X=19130 $Y=54570
X571 26 M11_M10_CDNS_7650684642119 $T=20090 63060 0 0 $X=19130 $Y=62780
X572 26 M11_M10_CDNS_7650684642119 $T=20090 73290 0 0 $X=19130 $Y=73010
X573 25 M11_M10_CDNS_7650684642119 $T=40560 14790 0 0 $X=39600 $Y=14510
X574 26 M11_M10_CDNS_7650684642119 $T=42240 37560 0 0 $X=41280 $Y=37280
X575 26 M11_M10_CDNS_7650684642119 $T=42240 46080 0 0 $X=41280 $Y=45800
X576 26 M11_M10_CDNS_7650684642119 $T=42240 54850 0 0 $X=41280 $Y=54570
X577 26 M11_M10_CDNS_7650684642119 $T=42240 63890 0 0 $X=41280 $Y=63610
X578 26 M11_M10_CDNS_7650684642119 $T=42240 83140 0 0 $X=41280 $Y=82860
X579 26 M11_M10_CDNS_7650684642119 $T=67370 29860 0 0 $X=66410 $Y=29580
X580 26 M11_M10_CDNS_7650684642119 $T=67370 37290 0 0 $X=66410 $Y=37010
X581 26 M11_M10_CDNS_7650684642119 $T=67370 46520 0 0 $X=66410 $Y=46240
X582 26 M11_M10_CDNS_7650684642119 $T=69160 53660 0 0 $X=68200 $Y=53380
X583 27 M11_M10_CDNS_7650684642119 $T=91890 5340 0 0 $X=90930 $Y=5060
X584 19 26 21 25 3 108 52 and2 $T=5890 68510 0 0 $X=3220 $Y=65930
X585 20 26 21 25 4 109 53 and2 $T=5890 78310 0 0 $X=3220 $Y=75730
X586 1 26 21 25 5 110 54 and2 $T=6190 47780 0 0 $X=3520 $Y=45200
X587 2 26 21 25 6 111 55 and2 $T=6190 57250 0 0 $X=3520 $Y=54670
X588 1 26 22 25 7 112 56 and2 $T=14410 42150 0 0 $X=11740 $Y=39570
X589 2 26 22 25 10 113 57 and2 $T=14510 52400 0 0 $X=11840 $Y=49820
X590 19 26 22 25 8 114 58 and2 $T=14510 61650 0 0 $X=11840 $Y=59070
X591 20 26 22 25 9 115 59 and2 $T=14510 71470 0 0 $X=11840 $Y=68890
X592 1 26 23 25 11 116 60 and2 $T=36030 34540 0 0 $X=33360 $Y=31960
X593 2 26 23 25 12 117 61 and2 $T=36880 43180 0 0 $X=34210 $Y=40600
X594 19 26 23 25 13 118 62 and2 $T=38080 51300 0 0 $X=35410 $Y=48720
X595 20 26 23 25 14 119 63 and2 $T=39970 59490 0 0 $X=37300 $Y=56910
X596 1 26 24 25 15 120 64 and2 $T=62470 24950 0 0 $X=59800 $Y=22370
X597 2 26 24 25 16 121 65 and2 $T=62710 34210 0 0 $X=60040 $Y=31630
X598 19 26 24 25 17 122 66 and2 $T=63260 42310 0 0 $X=60590 $Y=39730
X599 20 26 24 25 18 123 67 and2 $T=64690 50370 0 0 $X=62020 $Y=47790
X600 38 7 25 26 29 39 68 half_adder $T=19950 40210 0 0 $X=22250 $Y=40490
X601 9 3 25 26 28 37 70 half_adder $T=20250 64650 0 0 $X=22550 $Y=64930
X602 14 31 25 26 35 41 72 half_adder $T=45360 56090 0 0 $X=47660 $Y=56370
X603 18 34 25 26 47 44 74 half_adder $T=69570 48090 0 0 $X=71870 $Y=48370
X604 10 5 36 26 25 30 38 78 77 79
+ 76 full_adder $T=18880 47880 0 0 $X=20660 $Y=49130
X605 8 6 37 26 25 31 36 82 81 83
+ 80 full_adder $T=18880 56220 0 0 $X=20660 $Y=57470
X606 12 29 40 26 25 33 42 86 85 87
+ 84 full_adder $T=43990 39660 0 0 $X=45770 $Y=40910
X607 13 30 41 26 25 34 40 90 89 91
+ 88 full_adder $T=43990 47880 0 0 $X=45770 $Y=49130
X608 11 39 42 26 25 32 43 94 93 95
+ 92 full_adder $T=44590 31440 0 0 $X=46370 $Y=32690
X609 17 33 44 26 25 48 46 98 97 99
+ 96 full_adder $T=69190 39320 0 0 $X=70970 $Y=40570
X610 16 32 46 26 25 49 45 102 101 103
+ 100 full_adder $T=69850 30860 0 0 $X=71630 $Y=32110
X611 15 43 45 26 25 50 51 106 105 107
+ 104 full_adder $T=69860 22410 0 0 $X=71640 $Y=23660
M0 52 19 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3640 $Y=69440 $dt=1
M1 53 20 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3640 $Y=79240 $dt=1
M2 54 1 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3940 $Y=48710 $dt=1
M3 55 2 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3940 $Y=58180 $dt=1
M4 26 19 52 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4050 $Y=69440 $dt=1
M5 26 20 53 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4050 $Y=79240 $dt=1
M6 26 1 54 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4350 $Y=48710 $dt=1
M7 26 2 55 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=4350 $Y=58180 $dt=1
M8 52 21 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4940 $Y=69440 $dt=1
M9 53 21 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4940 $Y=79240 $dt=1
M10 54 21 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=5240 $Y=48710 $dt=1
M11 55 21 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=5240 $Y=58180 $dt=1
M12 56 1 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12160 $Y=43080 $dt=1
M13 57 2 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=53330 $dt=1
M14 58 19 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=62580 $dt=1
M15 59 20 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12260 $Y=72400 $dt=1
M16 26 1 56 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12570 $Y=43080 $dt=1
M17 26 2 57 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=53330 $dt=1
M18 26 19 58 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=62580 $dt=1
M19 26 20 59 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12670 $Y=72400 $dt=1
M20 56 22 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13460 $Y=43080 $dt=1
M21 57 22 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=53330 $dt=1
M22 58 22 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=62580 $dt=1
M23 59 22 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=13560 $Y=72400 $dt=1
M24 60 1 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=33780 $Y=35470 $dt=1
M25 26 1 60 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=34190 $Y=35470 $dt=1
M26 61 2 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=34630 $Y=44110 $dt=1
M27 26 2 61 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=35040 $Y=44110 $dt=1
M28 60 23 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=35080 $Y=35470 $dt=1
M29 62 19 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=35830 $Y=52230 $dt=1
M30 61 23 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=35930 $Y=44110 $dt=1
M31 26 19 62 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=36240 $Y=52230 $dt=1
M32 62 23 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=37130 $Y=52230 $dt=1
M33 63 20 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=37720 $Y=60420 $dt=1
M34 26 20 63 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=38130 $Y=60420 $dt=1
M35 63 23 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=39020 $Y=60420 $dt=1
M36 64 1 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=60220 $Y=25880 $dt=1
M37 65 2 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=60460 $Y=35140 $dt=1
M38 26 1 64 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=60630 $Y=25880 $dt=1
M39 26 2 65 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=60870 $Y=35140 $dt=1
M40 66 19 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=61010 $Y=43240 $dt=1
M41 26 19 66 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=61420 $Y=43240 $dt=1
M42 64 24 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=61520 $Y=25880 $dt=1
M43 65 24 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=61760 $Y=35140 $dt=1
M44 66 24 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=62310 $Y=43240 $dt=1
M45 67 20 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=62440 $Y=51300 $dt=1
M46 26 20 67 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=62850 $Y=51300 $dt=1
M47 67 24 26 26 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=63740 $Y=51300 $dt=1
.ends mult_auto
