* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : xor_auto                                     *
* Netlisted  : Thu Dec  4 09:31:52 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764862305972                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764862305972 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764862305972

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764862305973                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764862305973 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764862305973

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764862305974                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764862305974 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764862305974

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764862305975                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764862305975 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764862305975

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764862305970                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764862305970 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764862305970

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764862305971                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764862305971 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_764862305971

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
** N=4 EP=4 FDC=4
X0 2 3 1 2 2 nmos1v_CDNS_764862305970 $T=-60 -1520 0 0 $X=-480 $Y=-1720
X1 4 3 1 4 2 4 pmos1v_CDNS_764862305971 $T=-60 630 0 0 $X=-480 $Y=430
M0 3 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-60 $Y=630 $dt=1
M1 4 1 3 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=630 $dt=1
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor_auto                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor_auto 3 1 2 4 6 5
** N=6 EP=6 FDC=12
X0 1 M1_PO_CDNS_764862305972 $T=4460 3910 0 0 $X=4360 $Y=3790
X1 1 M1_PO_CDNS_764862305972 $T=4460 5790 0 0 $X=4360 $Y=5670
X2 2 M1_PO_CDNS_764862305972 $T=4870 1760 0 0 $X=4770 $Y=1640
X3 1 M1_PO_CDNS_764862305972 $T=4870 5790 0 0 $X=4770 $Y=5670
X4 3 M1_PO_CDNS_764862305972 $T=5760 2920 0 0 $X=5660 $Y=2800
X5 3 M2_M1_CDNS_764862305973 $T=4880 3450 0 0 $X=4750 $Y=3320
X6 4 M2_M1_CDNS_764862305973 $T=6240 3710 0 0 $X=6110 $Y=3580
X7 3 M2_M1_CDNS_764862305974 $T=4610 2640 0 0 $X=4480 $Y=2510
X8 3 M2_M1_CDNS_764862305974 $T=4660 4280 0 0 $X=4530 $Y=4150
X9 4 M2_M1_CDNS_764862305975 $T=4250 2340 0 0 $X=4170 $Y=2090
X10 4 M2_M1_CDNS_764862305975 $T=4250 4850 0 0 $X=4170 $Y=4600
X11 4 M2_M1_CDNS_764862305975 $T=5070 2340 0 0 $X=4990 $Y=2090
X12 4 M2_M1_CDNS_764862305975 $T=5070 4850 0 0 $X=4990 $Y=4600
X13 4 M2_M1_CDNS_764862305975 $T=5960 2340 0 0 $X=5880 $Y=2090
X14 4 M2_M1_CDNS_764862305975 $T=5960 4850 0 0 $X=5880 $Y=4600
X15 4 3 2 4 5 nmos1v_CDNS_764862305970 $T=4410 1980 0 0 $X=3990 $Y=1780
X16 2 4 3 2 5 nmos1v_CDNS_764862305970 $T=5710 1980 0 0 $X=5290 $Y=1780
X17 4 3 1 4 5 6 pmos1v_CDNS_764862305971 $T=4410 4130 0 0 $X=3990 $Y=3930
X18 1 4 3 1 5 6 pmos1v_CDNS_764862305971 $T=5710 4130 0 0 $X=5290 $Y=3930
X19 1 5 2 6 inv $T=3170 3500 0 0 $X=2690 $Y=1340
M0 3 1 4 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4410 $Y=4130 $dt=1
M1 4 1 3 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4820 $Y=4130 $dt=1
M2 4 3 1 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=5710 $Y=4130 $dt=1
M3 1 3 4 6 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=6120 $Y=4130 $dt=1
.ends xor_auto
