* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : and2                                         *
* Netlisted  : Sun Nov 30 13:51:59 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764532313970                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764532313970 S_source_0 D_drain_1 3 4 S_source_2 D_drain_3 B
** N=8 EP=7 FDC=3
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=37.8404 scb=0.0398877 scc=0.00354229 $X=0 $Y=0 $dt=1
M1 S_source_2 4 D_drain_1 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=32.9533 scb=0.0318315 scc=0.00282058 $X=410 $Y=0 $dt=1
M2 D_drain_3 D_drain_1 S_source_2 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=42.0058 scb=0.0446271 scc=0.00440038 $X=820 $Y=0 $dt=1
.ends pmos1v_CDNS_764532313970

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764532313971                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764532313971 S_source_0 D_drain_1 3 4 S_source_2 D_drain_3
** N=6 EP=6 FDC=3
M0 D_drain_1 3 S_source_0 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 S_source_2 4 D_drain_1 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 D_drain_3 S_source_0 S_source_2 S_source_2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
.ends nmos1v_CDNS_764532313971

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 A B OUT VDD VSS
** N=7 EP=5 FDC=6
X31 VDD 3 A B VDD OUT VDD pmos1v_CDNS_764532313970 $T=-460 820 0 0 $X=-880 $Y=620
X32 3 7 A B VSS OUT nmos1v_CDNS_764532313971 $T=-460 -1890 0 0 $X=-880 $Y=-2090
.ends and2
