* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : nand2_auto                                   *
* Netlisted  : Wed Dec  3 19:40:02 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764812396650                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764812396650 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764812396650

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764812396651                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764812396651 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764812396651

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764812396650                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764812396650 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_764812396650

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764812396651                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764812396651 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764812396651

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand2_auto                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand2_auto 1 2 4 5 6
** N=6 EP=5 FDC=8
X0 1 M1_PO_CDNS_764812396650 $T=2240 3700 0 0 $X=2140 $Y=3340
X1 2 M1_PO_CDNS_764812396650 $T=3540 3400 0 0 $X=3440 $Y=3040
X2 3 M2_M1_CDNS_764812396651 $T=2180 2120 0 0 $X=2100 $Y=1870
X3 4 M2_M1_CDNS_764812396651 $T=2590 4990 0 0 $X=2510 $Y=4740
X4 3 M2_M1_CDNS_764812396651 $T=3000 2120 0 0 $X=2920 $Y=1870
X5 3 M2_M1_CDNS_764812396651 $T=3480 2120 0 0 $X=3400 $Y=1870
X6 4 M2_M1_CDNS_764812396651 $T=3890 4990 0 0 $X=3810 $Y=4740
X7 3 M2_M1_CDNS_764812396651 $T=4300 2120 0 0 $X=4220 $Y=1870
X8 4 5 5 1 6 5 pmos1v_CDNS_764812396650 $T=2340 4270 0 0 $X=1920 $Y=4070
X9 4 5 5 2 6 5 pmos1v_CDNS_764812396650 $T=3640 4270 0 0 $X=3220 $Y=4070
X10 3 3 4 1 6 nmos1v_CDNS_764812396651 $T=2340 1400 0 0 $X=1920 $Y=1200
X11 3 3 6 2 6 nmos1v_CDNS_764812396651 $T=3640 1400 0 0 $X=3220 $Y=1200
M0 4 1 5 5 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2340 $Y=4270 $dt=1
M1 5 1 4 5 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.4011 scb=0.0195321 scc=0.00239618 $X=2750 $Y=4270 $dt=1
M2 4 2 5 5 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.4011 scb=0.0195321 scc=0.00239618 $X=3640 $Y=4270 $dt=1
M3 5 2 4 5 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=4050 $Y=4270 $dt=1
.ends nand2_auto
