* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mult                                         *
* Netlisted  : Sun Dec  7 18:49:31 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765154963930                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765154963930 S_source_0 S_source_2 D_drain_1 4 5
** N=5 EP=5 FDC=2
M0 D_drain_1 4 S_source_0 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 S_source_2 4 D_drain_1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765154963930

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765154963932                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765154963932 S_source_0 D_drain_1 3 S_source_2 5
** N=5 EP=5 FDC=2
M0 D_drain_1 3 S_source_0 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 S_source_2 3 D_drain_1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765154963932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv IN VDD OUT VSS
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X4 VSS OUT IN VSS VSS nmos1v_CDNS_765154963932 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 A VDD B VSS OUT 7
*.DEVICECLIMB
** N=7 EP=6 FDC=9
X10 6 6 7 A VSS nmos1v_CDNS_765154963930 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 6 6 VSS B VSS nmos1v_CDNS_765154963930 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X14 7 VDD OUT VSS inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 VDD B 7 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M1 OUT 7 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M2 VDD 7 OUT VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor B VDD VSS B_bar OUT A
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X8 OUT A B_bar OUT VSS nmos1v_CDNS_765154963932 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X9 B_bar OUT A B_bar VSS nmos1v_CDNS_765154963932 $T=800 -1920 0 0 $X=380 $Y=-2120
X10 B VDD B_bar VSS inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
M0 OUT B A VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 OUT A B VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 B A OUT VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765154963933                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765154963933 S_source_0 D_drain_1 3 S_source_2 D_drain_3 6 7 S_source_4 9
** N=9 EP=9 FDC=4
M0 D_drain_1 3 S_source_0 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 S_source_2 6 D_drain_1 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 D_drain_3 7 S_source_2 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 S_source_4 9 D_drain_3 S_source_2 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_765154963933

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765154963934                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765154963934 S_source_0 D_drain_1 S_source_2 4 5 D_drain_3 S_source_4 8 9 B
** N=11 EP=10 FDC=4
M0 D_drain_1 4 S_source_0 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 S_source_2 5 D_drain_1 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 D_drain_3 8 S_source_2 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 S_source_4 9 D_drain_3 B g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_765154963934

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network OUT P Ci VDD VSS P_bar A
** N=11 EP=7 FDC=8
X12 OUT 8 Ci VSS 9 P P_bar OUT A nmos1v_CDNS_765154963933 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 OUT 10 VDD Ci P_bar 11 OUT P A VDD pmos1v_CDNS_765154963934 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder B A Ci VDD VSS S Co
** N=15 EP=7 FDC=36
X14 10 VDD Co VSS inv $T=12350 3410 0 0 $X=11870 $Y=1250
X21 B VDD VSS 11 9 A xor $T=4170 3810 0 0 $X=1950 $Y=1250
X22 9 VDD VSS 8 S Ci xor $T=8070 3810 0 0 $X=5850 $Y=1250
X23 10 9 Ci VDD VSS 8 A fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 11 B VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 VDD B 11 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 A B 9 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 8 9 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 VDD 9 8 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 Ci 9 S VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 Co 10 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 VDD 10 Co VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder B A VSS VDD S Co
** N=9 EP=6 FDC=24
X6 A VDD B VSS Co 8 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X10 B VDD VSS 7 S A xor $T=4660 3560 0 0 $X=2440 $Y=1000
M0 7 B VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2860 $Y=3790 $dt=1
M1 VDD B 7 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3270 $Y=3790 $dt=1
M2 A B S VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4160 $Y=3790 $dt=1
M3 8 A VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6760 $Y=3790 $dt=1
M4 VDD A 8 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7170 $Y=3790 $dt=1
M5 8 B VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8060 $Y=3790 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mult                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mult A0 A1 A2 A3 B0 B1 B2 B3 P0 P1
+ P2 P3 P4 P5 P6 P7 VDD VSS
** N=143 EP=18 FDC=576
X584 A1 VDD B0 VSS 22 52 and2 $T=-8180 57870 0 0 $X=-10850 $Y=55290
X585 A0 VDD B0 VSS P0 53 and2 $T=-8180 67670 0 0 $X=-10850 $Y=65090
X586 A3 VDD B0 VSS 17 54 and2 $T=-7880 37140 0 0 $X=-10550 $Y=34560
X587 A2 VDD B0 VSS 18 55 and2 $T=-7880 46610 0 0 $X=-10550 $Y=44030
X588 A3 VDD B1 VSS 13 56 and2 $T=340 31510 0 0 $X=-2330 $Y=28930
X589 A2 VDD B1 VSS 16 57 and2 $T=440 41760 0 0 $X=-2230 $Y=39180
X590 A1 VDD B1 VSS 19 58 and2 $T=440 51010 0 0 $X=-2230 $Y=48430
X591 A0 VDD B1 VSS 21 59 and2 $T=440 60830 0 0 $X=-2230 $Y=58250
X592 A3 VDD B2 VSS 24 60 and2 $T=21960 23900 0 0 $X=19290 $Y=21320
X593 A2 VDD B2 VSS 23 61 and2 $T=22810 32540 0 0 $X=20140 $Y=29960
X594 A1 VDD B2 VSS 26 62 and2 $T=24010 40660 0 0 $X=21340 $Y=38080
X595 A0 VDD B2 VSS 27 63 and2 $T=25900 48850 0 0 $X=23230 $Y=46270
X596 A3 VDD B3 VSS 32 64 and2 $T=48400 14310 0 0 $X=45730 $Y=11730
X597 A2 VDD B3 VSS 31 65 and2 $T=48640 23570 0 0 $X=45970 $Y=20990
X598 A1 VDD B3 VSS 33 66 and2 $T=49190 31670 0 0 $X=46520 $Y=29090
X599 A0 VDD B3 VSS 35 67 and2 $T=50620 39730 0 0 $X=47950 $Y=37150
X600 16 17 14 VDD VSS 41 20 full_adder $T=4810 37240 0 0 $X=6590 $Y=38490
X601 19 18 15 VDD VSS 42 14 full_adder $T=4810 45580 0 0 $X=6590 $Y=46830
X602 23 40 28 VDD VSS 44 30 full_adder $T=29920 29020 0 0 $X=31700 $Y=30270
X603 26 41 29 VDD VSS 45 28 full_adder $T=29920 37240 0 0 $X=31700 $Y=38490
X604 24 25 30 VDD VSS 43 34 full_adder $T=30520 20800 0 0 $X=32300 $Y=22050
X605 33 44 36 VDD VSS P4 38 full_adder $T=55120 28680 0 0 $X=56900 $Y=29930
X606 31 43 38 VDD VSS P5 37 full_adder $T=55780 20220 0 0 $X=57560 $Y=21470
X607 32 34 37 VDD VSS P6 P7 full_adder $T=55790 11770 0 0 $X=57570 $Y=13020
X608 20 13 VSS VDD 40 25 half_adder $T=5880 29570 0 0 $X=8180 $Y=29850
X609 21 22 VSS VDD P1 15 half_adder $T=6180 54010 0 0 $X=8480 $Y=54290
X610 27 42 VSS VDD P2 29 half_adder $T=31290 45450 0 0 $X=33590 $Y=45730
X611 35 45 VSS VDD P3 36 half_adder $T=55500 37450 0 0 $X=57800 $Y=37730
M0 52 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10430 $Y=58800 $dt=1
M1 53 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10430 $Y=68600 $dt=1
M2 54 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10130 $Y=38070 $dt=1
M3 55 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10130 $Y=47540 $dt=1
M4 VDD A1 52 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-10020 $Y=58800 $dt=1
M5 VDD A0 53 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-10020 $Y=68600 $dt=1
M6 VDD A3 54 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-9720 $Y=38070 $dt=1
M7 VDD A2 55 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-9720 $Y=47540 $dt=1
M8 52 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-9130 $Y=58800 $dt=1
M9 53 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-9130 $Y=68600 $dt=1
M10 54 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-8830 $Y=38070 $dt=1
M11 55 B0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-8830 $Y=47540 $dt=1
M12 56 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1910 $Y=32440 $dt=1
M13 57 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1810 $Y=42690 $dt=1
M14 58 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1810 $Y=51940 $dt=1
M15 59 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1810 $Y=61760 $dt=1
M16 VDD A3 56 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1500 $Y=32440 $dt=1
M17 VDD A2 57 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1400 $Y=42690 $dt=1
M18 VDD A1 58 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1400 $Y=51940 $dt=1
M19 VDD A0 59 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1400 $Y=61760 $dt=1
M20 56 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-610 $Y=32440 $dt=1
M21 57 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-510 $Y=42690 $dt=1
M22 58 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-510 $Y=51940 $dt=1
M23 59 B1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-510 $Y=61760 $dt=1
M24 60 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=19710 $Y=24830 $dt=1
M25 VDD A3 60 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=20120 $Y=24830 $dt=1
M26 61 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=20560 $Y=33470 $dt=1
M27 VDD A2 61 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=20970 $Y=33470 $dt=1
M28 60 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=21010 $Y=24830 $dt=1
M29 62 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=21760 $Y=41590 $dt=1
M30 61 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=21860 $Y=33470 $dt=1
M31 VDD A1 62 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=22170 $Y=41590 $dt=1
M32 62 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=23060 $Y=41590 $dt=1
M33 63 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=23650 $Y=49780 $dt=1
M34 VDD A0 63 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=24060 $Y=49780 $dt=1
M35 63 B2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=24950 $Y=49780 $dt=1
M36 64 A3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=46150 $Y=15240 $dt=1
M37 65 A2 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=46390 $Y=24500 $dt=1
M38 VDD A3 64 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=46560 $Y=15240 $dt=1
M39 VDD A2 65 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=46800 $Y=24500 $dt=1
M40 66 A1 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=46940 $Y=32600 $dt=1
M41 VDD A1 66 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=47350 $Y=32600 $dt=1
M42 64 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=47450 $Y=15240 $dt=1
M43 65 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=47690 $Y=24500 $dt=1
M44 66 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=48240 $Y=32600 $dt=1
M45 67 A0 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=48370 $Y=40660 $dt=1
M46 VDD A0 67 VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=48780 $Y=40660 $dt=1
M47 67 B3 VDD VDD g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=49670 $Y=40660 $dt=1
.ends mult
