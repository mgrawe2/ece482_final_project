* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : c2mos                                        *
* Netlisted  : Sun Dec  7 19:23:32 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765157006931                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765157006931 S_source_0 2 D_drain_1 4
** N=4 EP=4 FDC=1
M0 D_drain_1 2 S_source_0 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765157006931

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765157006932                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765157006932 S_source_0 D_drain_1 3
** N=3 EP=3 FDC=1
M0 D_drain_1 3 S_source_0 D_drain_1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765157006932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: c2mos                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt c2mos CLK D Q RST VDD VSS
** N=12 EP=6 FDC=11
X21 VSS CLK 2 VSS nmos1v_CDNS_765157006931 $T=750 650 0 0 $X=330 $Y=450
X22 VSS D 11 VSS nmos1v_CDNS_765157006931 $T=2240 650 0 0 $X=1820 $Y=450
X23 11 2 3 VSS nmos1v_CDNS_765157006931 $T=3750 650 0 0 $X=3330 $Y=450
X24 VSS 3 12 VSS nmos1v_CDNS_765157006931 $T=5230 650 0 0 $X=4810 $Y=450
X25 12 CLK Q VSS nmos1v_CDNS_765157006931 $T=6720 650 0 0 $X=6300 $Y=450
X26 Q VSS RST nmos1v_CDNS_765157006932 $T=8210 170 0 0 $X=7790 $Y=-30
M0 2 CLK VDD VDD g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.27 scb=0.0231774 scc=0.00199917 $X=750 $Y=2360 $dt=1
M1 8 D VDD VDD g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=2240 $Y=2360 $dt=1
M2 3 CLK 8 VDD g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.7063 scb=0.016025 scc=0.00198503 $X=3740 $Y=2350 $dt=1
M3 9 3 VDD VDD g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=5230 $Y=2360 $dt=1
M4 Q 2 9 VDD g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.6749 scb=0.0214174 scc=0.0021813 $X=6720 $Y=2340 $dt=1
.ends c2mos
