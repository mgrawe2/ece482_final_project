* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : half_adder                                   *
* Netlisted  : Sun Nov 30 14:03:59 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764533033910                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764533033910 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764533033910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764533033911                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764533033911 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764533033911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764533033912                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764533033912 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764533033912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764533033913                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764533033913 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764533033913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764533033914                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764533033914 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764533033914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764533033915                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764533033915 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764533033915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764533033910                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764533033910 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.9282 scb=0.0134361 scc=0.000622896 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764533033910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764533033911                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764533033911 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=36.6317 scb=0.035909 scc=0.00335548 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764533033911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
** N=4 EP=4 FDC=2
X0 4 3 2 nmos1v_CDNS_764533033910 $T=-50 -540 0 0 $X=-470 $Y=-740
X1 1 3 2 4 1 pmos1v_CDNS_764533033911 $T=-50 460 0 0 $X=-470 $Y=260
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764533033912                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764533033912 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=0 $Y=0 $dt=1
M1 3 1 2 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=42.457 scb=0.04208 scc=0.00527302 $X=410 $Y=0 $dt=1
.ends pmos1v_CDNS_764533033912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764533033913                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764533033913 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=0 $Y=0 $dt=0
M1 3 1 2 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=5.15732 scb=0.00107852 scc=1.63215e-06 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764533033913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
** N=6 EP=6 FDC=6
X0 5 M2_M1_CDNS_764533033910 $T=360 650 0 0 $X=280 $Y=240
X1 5 M2_M1_CDNS_764533033910 $T=1260 650 0 0 $X=1180 $Y=240
X2 4 M1_PO_CDNS_764533033915 $T=850 -1090 0 0 $X=750 $Y=-1450
X3 3 M1_PO_CDNS_764533033915 $T=850 2390 0 0 $X=750 $Y=2030
X4 5 M1_PO_CDNS_764533033915 $T=1260 650 0 0 $X=1160 $Y=290
X5 1 3 4 2 inv $T=-790 -50 0 0 $X=-1590 $Y=-1230
X6 5 6 3 2 1 pmos1v_CDNS_764533033912 $T=660 1350 0 0 $X=240 $Y=1150
X7 5 6 4 2 nmos1v_CDNS_764533033913 $T=660 -340 0 0 $X=240 $Y=-540
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7645330339111                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7645330339111 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7645330339111

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7645330339112                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7645330339112 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7645330339112

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7645330339113                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7645330339113 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7645330339113

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7645330339114                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7645330339114 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7645330339114

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7645330339115                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7645330339115 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7645330339115

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_7645330339116                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_7645330339116 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_7645330339116

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_7645330339117                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_7645330339117 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_7645330339117

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_7645330339118                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_7645330339118 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_7645330339118

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_7645330339119                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_7645330339119 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_7645330339119

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764533033914                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764533033914 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=3
M0 2 3 1 8 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=5.5e-07 sca=26.2992 scb=0.0240146 scc=0.00255754 $X=0 $Y=0 $dt=1
M1 5 4 2 8 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.84e-14 PD=8e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=3.45e-07 sca=28.7383 scb=0.0277231 scc=0.00260208 $X=410 $Y=0 $dt=1
M2 6 2 5 8 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=5.5e-07 sb=1.4e-07 sca=39.2498 scb=0.0428135 scc=0.00408073 $X=820 $Y=0 $dt=1
.ends pmos1v_CDNS_764533033914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764533033915                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764533033915 1 2 3 4 5 6
** N=6 EP=6 FDC=3
M0 2 3 1 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
M1 5 4 2 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=410 $Y=0 $dt=0
M2 6 1 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=820 $Y=0 $dt=0
.ends nmos1v_CDNS_764533033915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7
** N=7 EP=7 FDC=6
X0 4 M2_M1_CDNS_764533033910 $T=-1500 -4280 0 0 $X=-1580 $Y=-4690
X1 3 M2_M1_CDNS_764533033910 $T=-990 -4280 0 0 $X=-1070 $Y=-4690
X2 5 M2_M1_CDNS_764533033910 $T=990 2710 0 0 $X=910 $Y=2300
X3 1 M2_M1_CDNS_764533033911 $T=-640 2480 0 0 $X=-1000 $Y=2350
X4 2 M2_M1_CDNS_764533033911 $T=680 -3080 0 0 $X=320 $Y=-3210
X5 3 M2_M1_CDNS_764533033912 $T=-560 200 0 0 $X=-640 $Y=-70
X6 4 M2_M1_CDNS_764533033912 $T=-150 -970 0 0 $X=-230 $Y=-1240
X7 3 M3_M2_CDNS_764533033913 $T=-560 200 0 0 $X=-640 $Y=-70
X8 4 M3_M2_CDNS_764533033913 $T=-150 -970 0 0 $X=-230 $Y=-1240
X9 4 M3_M2_CDNS_764533033914 $T=-1500 -4280 0 0 $X=-1580 $Y=-4690
X10 3 M3_M2_CDNS_764533033914 $T=-990 -4280 0 0 $X=-1070 $Y=-4690
X11 5 M3_M2_CDNS_764533033914 $T=990 2710 0 0 $X=910 $Y=2300
X12 3 M1_PO_CDNS_764533033915 $T=-560 200 0 0 $X=-660 $Y=-160
X13 4 M1_PO_CDNS_764533033915 $T=-150 -970 0 0 $X=-250 $Y=-1330
X14 6 M1_PO_CDNS_764533033915 $T=260 -270 0 0 $X=160 $Y=-630
X15 1 M3_M2_CDNS_7645330339111 $T=-640 2480 0 0 $X=-1000 $Y=2350
X16 2 M3_M2_CDNS_7645330339111 $T=680 -3080 0 0 $X=320 $Y=-3210
X17 1 M4_M3_CDNS_7645330339112 $T=-640 2480 0 0 $X=-1000 $Y=2350
X18 2 M4_M3_CDNS_7645330339112 $T=680 -3080 0 0 $X=320 $Y=-3210
X19 1 M5_M4_CDNS_7645330339113 $T=-640 2480 0 0 $X=-1000 $Y=2350
X20 2 M5_M4_CDNS_7645330339113 $T=680 -3080 0 0 $X=320 $Y=-3210
X21 1 M6_M5_CDNS_7645330339114 $T=-640 2480 0 0 $X=-1000 $Y=2350
X22 2 M6_M5_CDNS_7645330339114 $T=680 -3080 0 0 $X=320 $Y=-3210
X23 1 M7_M6_CDNS_7645330339115 $T=-640 2480 0 0 $X=-1000 $Y=2350
X24 2 M7_M6_CDNS_7645330339115 $T=680 -3080 0 0 $X=320 $Y=-3210
X25 1 M8_M7_CDNS_7645330339116 $T=-640 2480 0 0 $X=-1000 $Y=2350
X26 2 M8_M7_CDNS_7645330339116 $T=680 -3080 0 0 $X=320 $Y=-3210
X27 1 M9_M8_CDNS_7645330339117 $T=-640 2480 0 0 $X=-1000 $Y=2350
X28 2 M9_M8_CDNS_7645330339117 $T=680 -3080 0 0 $X=320 $Y=-3210
X29 1 M10_M9_CDNS_7645330339118 $T=-630 2470 0 0 $X=-1590 $Y=2190
X30 2 M10_M9_CDNS_7645330339118 $T=700 -3080 0 0 $X=-260 $Y=-3360
X31 1 M11_M10_CDNS_7645330339119 $T=-630 2470 0 0 $X=-1590 $Y=2190
X32 2 M11_M10_CDNS_7645330339119 $T=700 -3080 0 0 $X=-260 $Y=-3360
X33 1 6 3 4 1 5 2 1 pmos1v_CDNS_764533033914 $T=-460 820 0 0 $X=-880 $Y=620
X34 6 7 3 4 2 5 nmos1v_CDNS_764533033915 $T=-460 -1890 0 0 $X=-880 $Y=-2090
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 2 1 7 3 4 5
** N=9 EP=6 FDC=12
X0 1 M2_M1_CDNS_764533033910 $T=-4170 -2510 0 0 $X=-4250 $Y=-2920
X1 1 M2_M1_CDNS_764533033910 $T=-4170 440 0 0 $X=-4250 $Y=30
X2 2 M2_M1_CDNS_764533033910 $T=-1860 -2510 0 0 $X=-1940 $Y=-2920
X3 3 M2_M1_CDNS_764533033910 $T=-1450 3410 0 0 $X=-1530 $Y=3000
X4 4 M2_M1_CDNS_764533033911 $T=-3220 1460 0 0 $X=-3580 $Y=1330
X5 4 M2_M1_CDNS_764533033911 $T=620 2430 0 0 $X=260 $Y=2300
X6 3 M2_M1_CDNS_764533033912 $T=-1450 460 0 0 $X=-1530 $Y=190
X7 3 M3_M2_CDNS_764533033913 $T=-1450 460 0 0 $X=-1530 $Y=190
X8 1 M3_M2_CDNS_764533033914 $T=-4170 -2510 0 0 $X=-4250 $Y=-2920
X9 2 M3_M2_CDNS_764533033914 $T=-1860 -2510 0 0 $X=-1940 $Y=-2920
X10 2 M3_M2_CDNS_764533033914 $T=-1860 720 0 0 $X=-1940 $Y=310
X11 3 M3_M2_CDNS_764533033914 $T=-1450 3410 0 0 $X=-1530 $Y=3000
X12 4 5 1 6 2 3 xor $T=-2220 70 0 0 $X=-4090 $Y=-1380
X13 4 5 2 1 7 8 9 and2 $T=630 630 0 0 $X=-960 $Y=-4060
.ends half_adder
