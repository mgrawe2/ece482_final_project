* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mult                                         *
* Netlisted  : Sun Dec  7 18:49:31 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_765154963930                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_765154963930 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_765154963930

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765154963931                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765154963931 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765154963931

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_765154963932                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_765154963932 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_765154963932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_765154963933                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_765154963933 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_765154963933

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_765154963934                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_765154963934 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_765154963934

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_765154963935                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_765154963935 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_765154963935

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_765154963936                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_765154963936 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_765154963936

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765154963937                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765154963937 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765154963937

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765154963938                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765154963938 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765154963938

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765154963939                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765154963939 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765154963939

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7651549639310                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7651549639310 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7651549639310

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651549639311                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651549639311 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651549639311

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651549639312                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651549639312 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651549639312

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651549639313                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651549639313 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651549639313

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651549639314                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651549639314 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651549639314

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651549639315                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651549639315 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651549639315

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651549639317                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651549639317 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651549639317

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651549639318                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651549639318 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651549639318

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651549639319                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651549639319 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651549639319

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_7651549639320                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_7651549639320 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_7651549639320

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651549639321                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651549639321 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651549639321

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_7651549639322                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_7651549639322 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_7651549639322

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651549639323                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651549639323 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651549639323

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765154963930                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765154963930 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765154963930

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765154963931                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765154963931 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_765154963931

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765154963932                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765154963932 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765154963932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X0 2 M1_NWELL_CDNS_7651549639320 $T=190 2570 0 0 $X=-230 $Y=2270
X1 4 M1_PSUB_CDNS_7651549639322 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 1 M1_PO_CDNS_7651549639323 $T=-160 30 0 0 $X=-260 $Y=-330
X3 2 3 1 2 4 2 pmos1v_CDNS_765154963931 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 3 1 4 4 nmos1v_CDNS_765154963932 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=9
X0 2 M1_NWELL_CDNS_7651549639320 $T=-1350 2870 0 0 $X=-1770 $Y=2570
X1 6 M2_M1_CDNS_7651549639321 $T=-2410 -1220 0 0 $X=-2490 $Y=-1470
X2 7 M2_M1_CDNS_7651549639321 $T=-2000 1650 0 0 $X=-2080 $Y=1400
X3 6 M2_M1_CDNS_7651549639321 $T=-1590 -1220 0 0 $X=-1670 $Y=-1470
X4 6 M2_M1_CDNS_7651549639321 $T=-1110 -1220 0 0 $X=-1190 $Y=-1470
X5 7 M2_M1_CDNS_7651549639321 $T=-700 1650 0 0 $X=-780 $Y=1400
X6 6 M2_M1_CDNS_7651549639321 $T=-290 -1220 0 0 $X=-370 $Y=-1470
X7 4 M1_PSUB_CDNS_7651549639322 $T=-700 -2440 0 0 $X=-1080 $Y=-2580
X8 1 M1_PO_CDNS_7651549639323 $T=-2350 360 0 0 $X=-2450 $Y=0
X9 3 M1_PO_CDNS_7651549639323 $T=-1050 60 0 0 $X=-1150 $Y=-300
X10 6 6 7 1 4 nmos1v_CDNS_765154963930 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 6 6 4 3 4 nmos1v_CDNS_765154963930 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X12 2 7 1 2 4 2 pmos1v_CDNS_765154963931 $T=-2250 930 0 0 $X=-2670 $Y=730
X13 2 7 3 2 4 2 pmos1v_CDNS_765154963931 $T=-950 930 0 0 $X=-1370 $Y=730
X14 7 2 5 4 inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 2 3 7 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M1 5 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M2 2 7 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651549639324                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651549639324 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651549639324

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651549639325                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651549639325 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651549639325

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651549639326                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651549639326 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651549639326

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651549639329                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651549639329 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651549639329

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X0 5 M2_M1_CDNS_7651549639321 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X1 5 M2_M1_CDNS_7651549639321 $T=-660 950 0 0 $X=-740 $Y=700
X2 5 M2_M1_CDNS_7651549639321 $T=160 -1560 0 0 $X=80 $Y=-1810
X3 5 M2_M1_CDNS_7651549639321 $T=160 950 0 0 $X=80 $Y=700
X4 5 M2_M1_CDNS_7651549639321 $T=1050 -1560 0 0 $X=970 $Y=-1810
X5 5 M2_M1_CDNS_7651549639321 $T=1050 950 0 0 $X=970 $Y=700
X6 5 6 1 5 3 2 pmos1v_CDNS_765154963931 $T=-500 230 0 0 $X=-920 $Y=30
X7 1 5 6 1 3 2 pmos1v_CDNS_765154963931 $T=800 230 0 0 $X=380 $Y=30
X8 5 6 4 5 3 nmos1v_CDNS_765154963932 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X9 4 5 6 4 3 nmos1v_CDNS_765154963932 $T=800 -1920 0 0 $X=380 $Y=-2120
X10 1 2 4 3 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
X11 6 M2_M1_CDNS_7651549639325 $T=-30 -450 0 0 $X=-160 $Y=-580
X12 5 M2_M1_CDNS_7651549639325 $T=1330 -190 0 0 $X=1200 $Y=-320
X13 6 M2_M1_CDNS_7651549639326 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X14 6 M2_M1_CDNS_7651549639326 $T=-250 380 0 0 $X=-380 $Y=250
X15 1 M1_PO_CDNS_7651549639329 $T=-450 10 0 0 $X=-550 $Y=-110
X16 1 M1_PO_CDNS_7651549639329 $T=-450 1890 0 0 $X=-550 $Y=1770
X17 4 M1_PO_CDNS_7651549639329 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X18 1 M1_PO_CDNS_7651549639329 $T=-40 1890 0 0 $X=-140 $Y=1770
X19 6 M1_PO_CDNS_7651549639329 $T=850 -980 0 0 $X=750 $Y=-1100
M0 5 1 6 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 5 6 1 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 1 6 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765154963933                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765154963933 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_765154963933

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765154963934                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765154963934 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_765154963934

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=8
X0 1 M2_M1_CDNS_7651549639315 $T=-830 -970 0 0 $X=-910 $Y=-1100
X1 2 M2_M1_CDNS_7651549639315 $T=-220 -60 0 0 $X=-300 $Y=-190
X2 2 M2_M1_CDNS_7651549639315 $T=200 730 0 0 $X=120 $Y=600
X3 1 M2_M1_CDNS_7651549639315 $T=810 -970 0 0 $X=730 $Y=-1100
X4 4 M1_NWELL_CDNS_7651549639320 $T=-10 2990 0 0 $X=-430 $Y=2690
X5 5 M1_PSUB_CDNS_7651549639322 $T=0 -1600 0 0 $X=-380 $Y=-1740
X6 3 M1_PO_CDNS_7651549639323 $T=-590 550 0 0 $X=-690 $Y=190
X7 7 M1_PO_CDNS_7651549639323 $T=570 550 0 0 $X=470 $Y=190
X8 2 M1_PO_CDNS_7651549639329 $T=-220 -60 0 0 $X=-320 $Y=-180
X9 6 M1_PO_CDNS_7651549639329 $T=-210 730 0 0 $X=-310 $Y=610
X10 6 M1_PO_CDNS_7651549639329 $T=190 -60 0 0 $X=90 $Y=-180
X11 2 M1_PO_CDNS_7651549639329 $T=200 730 0 0 $X=100 $Y=610
X12 1 8 3 5 9 2 6 1 7 nmos1v_CDNS_765154963933 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 1 10 4 3 6 11 1 2 7 5
+ 4 pmos1v_CDNS_765154963934 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 1 2 3 4 5 6 7 8 9 10
+ 11
** N=15 EP=11 FDC=36
X0 1 M3_M2_CDNS_7651549639314 $T=2270 3860 0 0 $X=2190 $Y=3730
X1 2 M3_M2_CDNS_7651549639314 $T=5790 3080 0 0 $X=5710 $Y=2950
X2 6 M3_M2_CDNS_7651549639314 $T=9120 4760 0 0 $X=9040 $Y=4630
X3 2 M3_M2_CDNS_7651549639314 $T=11410 2940 0 0 $X=11330 $Y=2810
X4 7 M3_M2_CDNS_7651549639314 $T=12920 3510 0 0 $X=12840 $Y=3380
X5 2 M2_M1_CDNS_7651549639315 $T=5250 3070 0 0 $X=5170 $Y=2940
X6 8 M2_M1_CDNS_7651549639315 $T=9530 2380 0 0 $X=9450 $Y=2250
X7 9 M2_M1_CDNS_7651549639315 $T=9530 5090 0 0 $X=9450 $Y=4960
X8 4 M2_M1_CDNS_7651549639315 $T=10820 5970 0 0 $X=10740 $Y=5840
X9 8 M2_M1_CDNS_7651549639315 $T=11040 2940 0 0 $X=10960 $Y=2810
X10 2 M2_M1_CDNS_7651549639315 $T=11390 3320 0 0 $X=11310 $Y=3190
X11 7 M2_M1_CDNS_7651549639315 $T=12920 3510 0 0 $X=12840 $Y=3380
X12 2 M4_M3_CDNS_7651549639319 $T=6980 3080 0 0 $X=6900 $Y=2950
X13 2 M4_M3_CDNS_7651549639319 $T=10140 2970 0 0 $X=10060 $Y=2840
X14 10 4 7 5 inv $T=12350 3410 0 0 $X=11870 $Y=1250
X15 3 M3_M2_CDNS_7651549639324 $T=7300 3360 0 0 $X=7170 $Y=3230
X16 3 M3_M2_CDNS_7651549639324 $T=10110 3640 0 0 $X=9980 $Y=3510
X17 4 M2_M1_CDNS_7651549639325 $T=6470 5920 0 0 $X=6340 $Y=5790
X18 3 M2_M1_CDNS_7651549639325 $T=7620 3360 0 0 $X=7490 $Y=3230
X19 3 M2_M1_CDNS_7651549639325 $T=10320 3640 0 0 $X=10190 $Y=3510
X20 4 M2_M1_CDNS_7651549639326 $T=3420 5920 0 0 $X=3290 $Y=5790
X21 1 4 5 11 9 2 xor $T=4170 3810 0 0 $X=1950 $Y=1250
X22 9 4 5 8 6 3 xor $T=8070 3810 0 0 $X=5850 $Y=1250
X23 10 9 3 4 5 8 2 12 13 14
+ 15 fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 11 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 4 1 11 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 2 1 9 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 8 9 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 4 9 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 3 9 6 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 7 10 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 4 10 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 7
** N=9 EP=7 FDC=24
X0 1 M3_M2_CDNS_7651549639314 $T=2760 3570 0 0 $X=2680 $Y=3440
X1 2 M3_M2_CDNS_7651549639314 $T=4630 3110 0 0 $X=4550 $Y=2980
X2 6 M3_M2_CDNS_7651549639314 $T=9970 3310 0 0 $X=9890 $Y=3180
X3 5 M3_M2_CDNS_7651549639314 $T=10180 2730 0 0 $X=10100 $Y=2600
X4 6 M2_M1_CDNS_7651549639315 $T=9970 3310 0 0 $X=9890 $Y=3180
X5 5 M2_M1_CDNS_7651549639315 $T=10180 2730 0 0 $X=10100 $Y=2600
X6 2 4 1 3 6 9 8 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X7 1 M2_M1_CDNS_7651549639325 $T=2760 2580 0 0 $X=2630 $Y=2450
X8 1 M2_M1_CDNS_7651549639325 $T=7960 2810 0 0 $X=7830 $Y=2680
X9 5 M2_M1_CDNS_7651549639326 $T=6360 3430 0 0 $X=6230 $Y=3300
X10 1 4 3 7 5 2 xor $T=4660 3560 0 0 $X=2440 $Y=1000
M0 7 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2860 $Y=3790 $dt=1
M1 4 1 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3270 $Y=3790 $dt=1
M2 2 1 5 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4160 $Y=3790 $dt=1
M3 8 2 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6760 $Y=3790 $dt=1
M4 4 2 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7170 $Y=3790 $dt=1
M5 8 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8060 $Y=3790 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mult                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mult 8 6 5 4 9 10 11 12 39 7
+ 46 51 47 48 49 50 1 2
** N=143 EP=18 FDC=576
X0 1 M11_M10_CDNS_765154963930 $T=-4370 38930 0 0 $X=-5330 $Y=38650
X1 1 M11_M10_CDNS_765154963930 $T=-4370 45380 0 0 $X=-5330 $Y=45100
X2 1 M11_M10_CDNS_765154963930 $T=-4370 60080 0 0 $X=-5330 $Y=59800
X3 1 M11_M10_CDNS_765154963930 $T=-3860 70340 0 0 $X=-4820 $Y=70060
X4 1 M11_M10_CDNS_765154963930 $T=6020 35670 0 0 $X=5060 $Y=35390
X5 1 M11_M10_CDNS_765154963930 $T=6020 44210 0 0 $X=5060 $Y=43930
X6 1 M11_M10_CDNS_765154963930 $T=6020 52420 0 0 $X=5060 $Y=52140
X7 1 M11_M10_CDNS_765154963930 $T=6020 62650 0 0 $X=5060 $Y=62370
X8 2 M11_M10_CDNS_765154963930 $T=26490 4150 0 0 $X=25530 $Y=3870
X9 1 M11_M10_CDNS_765154963930 $T=28170 26920 0 0 $X=27210 $Y=26640
X10 1 M11_M10_CDNS_765154963930 $T=28170 35440 0 0 $X=27210 $Y=35160
X11 1 M11_M10_CDNS_765154963930 $T=28170 44210 0 0 $X=27210 $Y=43930
X12 1 M11_M10_CDNS_765154963930 $T=28170 53250 0 0 $X=27210 $Y=52970
X13 1 M11_M10_CDNS_765154963930 $T=28170 72500 0 0 $X=27210 $Y=72220
X14 1 M11_M10_CDNS_765154963930 $T=53300 19220 0 0 $X=52340 $Y=18940
X15 1 M11_M10_CDNS_765154963930 $T=53300 26650 0 0 $X=52340 $Y=26370
X16 1 M11_M10_CDNS_765154963930 $T=53300 35880 0 0 $X=52340 $Y=35600
X17 1 M11_M10_CDNS_765154963930 $T=55090 43020 0 0 $X=54130 $Y=42740
X18 3 M11_M10_CDNS_765154963930 $T=77820 -5300 0 0 $X=76860 $Y=-5580
X19 2 M5_M4_CDNS_765154963931 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X20 2 M5_M4_CDNS_765154963931 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X21 2 M5_M4_CDNS_765154963931 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X22 2 M5_M4_CDNS_765154963931 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X23 1 M5_M4_CDNS_765154963931 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X24 1 M5_M4_CDNS_765154963931 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X25 1 M5_M4_CDNS_765154963931 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X26 1 M5_M4_CDNS_765154963931 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X27 2 M5_M4_CDNS_765154963931 $T=1340 28530 0 0 $X=980 $Y=28400
X28 2 M5_M4_CDNS_765154963931 $T=1340 38870 0 0 $X=980 $Y=38740
X29 2 M5_M4_CDNS_765154963931 $T=2350 48710 0 0 $X=1990 $Y=48580
X30 2 M5_M4_CDNS_765154963931 $T=2350 58460 0 0 $X=1990 $Y=58330
X31 1 M5_M4_CDNS_765154963931 $T=6020 35670 0 0 $X=5660 $Y=35540
X32 1 M5_M4_CDNS_765154963931 $T=6020 44210 0 0 $X=5660 $Y=44080
X33 1 M5_M4_CDNS_765154963931 $T=6020 52420 0 0 $X=5660 $Y=52290
X34 1 M5_M4_CDNS_765154963931 $T=6020 62650 0 0 $X=5660 $Y=62520
X35 2 M5_M4_CDNS_765154963931 $T=7810 29790 0 0 $X=7450 $Y=29660
X36 2 M5_M4_CDNS_765154963931 $T=7810 38630 0 0 $X=7450 $Y=38500
X37 2 M5_M4_CDNS_765154963931 $T=7810 45970 0 0 $X=7450 $Y=45840
X38 2 M5_M4_CDNS_765154963931 $T=7810 54500 0 0 $X=7450 $Y=54370
X39 2 M5_M4_CDNS_765154963931 $T=23540 29510 0 0 $X=23180 $Y=29380
X40 2 M5_M4_CDNS_765154963931 $T=23540 36860 0 0 $X=23180 $Y=36730
X41 2 M5_M4_CDNS_765154963931 $T=24360 21640 0 0 $X=24000 $Y=21510
X42 2 M5_M4_CDNS_765154963931 $T=26800 45560 0 0 $X=26440 $Y=45430
X43 1 M5_M4_CDNS_765154963931 $T=28170 26920 0 0 $X=27810 $Y=26790
X44 1 M5_M4_CDNS_765154963931 $T=28170 35440 0 0 $X=27810 $Y=35310
X45 1 M5_M4_CDNS_765154963931 $T=28170 44210 0 0 $X=27810 $Y=44080
X46 1 M5_M4_CDNS_765154963931 $T=28170 53250 0 0 $X=27810 $Y=53120
X47 1 M5_M4_CDNS_765154963931 $T=28170 72500 0 0 $X=27810 $Y=72370
X48 2 M5_M4_CDNS_765154963931 $T=30470 38630 0 0 $X=30110 $Y=38500
X49 2 M5_M4_CDNS_765154963931 $T=33760 21470 0 0 $X=33400 $Y=21340
X50 2 M5_M4_CDNS_765154963931 $T=33760 29680 0 0 $X=33400 $Y=29550
X51 2 M5_M4_CDNS_765154963931 $T=34980 45870 0 0 $X=34620 $Y=45740
X52 2 M5_M4_CDNS_765154963931 $T=50880 20850 0 0 $X=50520 $Y=20720
X53 2 M5_M4_CDNS_765154963931 $T=50880 28780 0 0 $X=50520 $Y=28650
X54 2 M5_M4_CDNS_765154963931 $T=50880 36650 0 0 $X=50520 $Y=36520
X55 2 M5_M4_CDNS_765154963931 $T=51050 12420 0 0 $X=50690 $Y=12290
X56 1 M5_M4_CDNS_765154963931 $T=53300 19220 0 0 $X=52940 $Y=19090
X57 1 M5_M4_CDNS_765154963931 $T=53300 26650 0 0 $X=52940 $Y=26520
X58 1 M5_M4_CDNS_765154963931 $T=53300 35880 0 0 $X=52940 $Y=35750
X59 1 M5_M4_CDNS_765154963931 $T=55090 43020 0 0 $X=54730 $Y=42890
X60 2 M5_M4_CDNS_765154963931 $T=57390 12420 0 0 $X=57030 $Y=12290
X61 2 M5_M4_CDNS_765154963931 $T=57390 20810 0 0 $X=57030 $Y=20680
X62 2 M5_M4_CDNS_765154963931 $T=57390 29200 0 0 $X=57030 $Y=29070
X63 2 M5_M4_CDNS_765154963931 $T=57390 37590 0 0 $X=57030 $Y=37460
X64 3 M5_M4_CDNS_765154963931 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X65 2 M6_M5_CDNS_765154963932 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X66 2 M6_M5_CDNS_765154963932 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X67 2 M6_M5_CDNS_765154963932 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X68 2 M6_M5_CDNS_765154963932 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X69 1 M6_M5_CDNS_765154963932 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X70 1 M6_M5_CDNS_765154963932 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X71 1 M6_M5_CDNS_765154963932 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X72 1 M6_M5_CDNS_765154963932 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X73 2 M6_M5_CDNS_765154963932 $T=1340 28530 0 0 $X=980 $Y=28400
X74 2 M6_M5_CDNS_765154963932 $T=1340 38870 0 0 $X=980 $Y=38740
X75 2 M6_M5_CDNS_765154963932 $T=2350 48710 0 0 $X=1990 $Y=48580
X76 2 M6_M5_CDNS_765154963932 $T=2350 58460 0 0 $X=1990 $Y=58330
X77 1 M6_M5_CDNS_765154963932 $T=6020 35670 0 0 $X=5660 $Y=35540
X78 1 M6_M5_CDNS_765154963932 $T=6020 44210 0 0 $X=5660 $Y=44080
X79 1 M6_M5_CDNS_765154963932 $T=6020 52420 0 0 $X=5660 $Y=52290
X80 1 M6_M5_CDNS_765154963932 $T=6020 62650 0 0 $X=5660 $Y=62520
X81 2 M6_M5_CDNS_765154963932 $T=7810 29790 0 0 $X=7450 $Y=29660
X82 2 M6_M5_CDNS_765154963932 $T=7810 38630 0 0 $X=7450 $Y=38500
X83 2 M6_M5_CDNS_765154963932 $T=7810 45970 0 0 $X=7450 $Y=45840
X84 2 M6_M5_CDNS_765154963932 $T=7810 54500 0 0 $X=7450 $Y=54370
X85 2 M6_M5_CDNS_765154963932 $T=23540 29510 0 0 $X=23180 $Y=29380
X86 2 M6_M5_CDNS_765154963932 $T=23540 36860 0 0 $X=23180 $Y=36730
X87 2 M6_M5_CDNS_765154963932 $T=24360 21640 0 0 $X=24000 $Y=21510
X88 2 M6_M5_CDNS_765154963932 $T=26800 45560 0 0 $X=26440 $Y=45430
X89 1 M6_M5_CDNS_765154963932 $T=28170 26920 0 0 $X=27810 $Y=26790
X90 1 M6_M5_CDNS_765154963932 $T=28170 35440 0 0 $X=27810 $Y=35310
X91 1 M6_M5_CDNS_765154963932 $T=28170 44210 0 0 $X=27810 $Y=44080
X92 1 M6_M5_CDNS_765154963932 $T=28170 53250 0 0 $X=27810 $Y=53120
X93 1 M6_M5_CDNS_765154963932 $T=28170 72500 0 0 $X=27810 $Y=72370
X94 2 M6_M5_CDNS_765154963932 $T=30470 38630 0 0 $X=30110 $Y=38500
X95 2 M6_M5_CDNS_765154963932 $T=33760 21470 0 0 $X=33400 $Y=21340
X96 2 M6_M5_CDNS_765154963932 $T=33760 29680 0 0 $X=33400 $Y=29550
X97 2 M6_M5_CDNS_765154963932 $T=34980 45870 0 0 $X=34620 $Y=45740
X98 2 M6_M5_CDNS_765154963932 $T=50880 20850 0 0 $X=50520 $Y=20720
X99 2 M6_M5_CDNS_765154963932 $T=50880 28780 0 0 $X=50520 $Y=28650
X100 2 M6_M5_CDNS_765154963932 $T=50880 36650 0 0 $X=50520 $Y=36520
X101 2 M6_M5_CDNS_765154963932 $T=51050 12420 0 0 $X=50690 $Y=12290
X102 1 M6_M5_CDNS_765154963932 $T=53300 19220 0 0 $X=52940 $Y=19090
X103 1 M6_M5_CDNS_765154963932 $T=53300 26650 0 0 $X=52940 $Y=26520
X104 1 M6_M5_CDNS_765154963932 $T=53300 35880 0 0 $X=52940 $Y=35750
X105 1 M6_M5_CDNS_765154963932 $T=55090 43020 0 0 $X=54730 $Y=42890
X106 2 M6_M5_CDNS_765154963932 $T=57390 12420 0 0 $X=57030 $Y=12290
X107 2 M6_M5_CDNS_765154963932 $T=57390 20810 0 0 $X=57030 $Y=20680
X108 2 M6_M5_CDNS_765154963932 $T=57390 29200 0 0 $X=57030 $Y=29070
X109 2 M6_M5_CDNS_765154963932 $T=57390 37590 0 0 $X=57030 $Y=37460
X110 3 M6_M5_CDNS_765154963932 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X111 2 M7_M6_CDNS_765154963933 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X112 2 M7_M6_CDNS_765154963933 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X113 2 M7_M6_CDNS_765154963933 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X114 2 M7_M6_CDNS_765154963933 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X115 1 M7_M6_CDNS_765154963933 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X116 1 M7_M6_CDNS_765154963933 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X117 1 M7_M6_CDNS_765154963933 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X118 1 M7_M6_CDNS_765154963933 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X119 2 M7_M6_CDNS_765154963933 $T=1340 28530 0 0 $X=980 $Y=28400
X120 2 M7_M6_CDNS_765154963933 $T=1340 38870 0 0 $X=980 $Y=38740
X121 2 M7_M6_CDNS_765154963933 $T=2350 48710 0 0 $X=1990 $Y=48580
X122 2 M7_M6_CDNS_765154963933 $T=2350 58460 0 0 $X=1990 $Y=58330
X123 1 M7_M6_CDNS_765154963933 $T=6020 35670 0 0 $X=5660 $Y=35540
X124 1 M7_M6_CDNS_765154963933 $T=6020 44210 0 0 $X=5660 $Y=44080
X125 1 M7_M6_CDNS_765154963933 $T=6020 52420 0 0 $X=5660 $Y=52290
X126 1 M7_M6_CDNS_765154963933 $T=6020 62650 0 0 $X=5660 $Y=62520
X127 2 M7_M6_CDNS_765154963933 $T=7810 29790 0 0 $X=7450 $Y=29660
X128 2 M7_M6_CDNS_765154963933 $T=7810 38630 0 0 $X=7450 $Y=38500
X129 2 M7_M6_CDNS_765154963933 $T=7810 45970 0 0 $X=7450 $Y=45840
X130 2 M7_M6_CDNS_765154963933 $T=7810 54500 0 0 $X=7450 $Y=54370
X131 2 M7_M6_CDNS_765154963933 $T=23540 29510 0 0 $X=23180 $Y=29380
X132 2 M7_M6_CDNS_765154963933 $T=23540 36860 0 0 $X=23180 $Y=36730
X133 2 M7_M6_CDNS_765154963933 $T=24360 21640 0 0 $X=24000 $Y=21510
X134 2 M7_M6_CDNS_765154963933 $T=26800 45560 0 0 $X=26440 $Y=45430
X135 1 M7_M6_CDNS_765154963933 $T=28170 26920 0 0 $X=27810 $Y=26790
X136 1 M7_M6_CDNS_765154963933 $T=28170 35440 0 0 $X=27810 $Y=35310
X137 1 M7_M6_CDNS_765154963933 $T=28170 44210 0 0 $X=27810 $Y=44080
X138 1 M7_M6_CDNS_765154963933 $T=28170 53250 0 0 $X=27810 $Y=53120
X139 1 M7_M6_CDNS_765154963933 $T=28170 72500 0 0 $X=27810 $Y=72370
X140 2 M7_M6_CDNS_765154963933 $T=30470 38630 0 0 $X=30110 $Y=38500
X141 2 M7_M6_CDNS_765154963933 $T=33760 21470 0 0 $X=33400 $Y=21340
X142 2 M7_M6_CDNS_765154963933 $T=33760 29680 0 0 $X=33400 $Y=29550
X143 2 M7_M6_CDNS_765154963933 $T=34980 45870 0 0 $X=34620 $Y=45740
X144 2 M7_M6_CDNS_765154963933 $T=50880 20850 0 0 $X=50520 $Y=20720
X145 2 M7_M6_CDNS_765154963933 $T=50880 28780 0 0 $X=50520 $Y=28650
X146 2 M7_M6_CDNS_765154963933 $T=50880 36650 0 0 $X=50520 $Y=36520
X147 2 M7_M6_CDNS_765154963933 $T=51050 12420 0 0 $X=50690 $Y=12290
X148 1 M7_M6_CDNS_765154963933 $T=53300 19220 0 0 $X=52940 $Y=19090
X149 1 M7_M6_CDNS_765154963933 $T=53300 26650 0 0 $X=52940 $Y=26520
X150 1 M7_M6_CDNS_765154963933 $T=53300 35880 0 0 $X=52940 $Y=35750
X151 1 M7_M6_CDNS_765154963933 $T=55090 43020 0 0 $X=54730 $Y=42890
X152 2 M7_M6_CDNS_765154963933 $T=57390 12420 0 0 $X=57030 $Y=12290
X153 2 M7_M6_CDNS_765154963933 $T=57390 20810 0 0 $X=57030 $Y=20680
X154 2 M7_M6_CDNS_765154963933 $T=57390 29200 0 0 $X=57030 $Y=29070
X155 2 M7_M6_CDNS_765154963933 $T=57390 37590 0 0 $X=57030 $Y=37460
X156 3 M7_M6_CDNS_765154963933 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X157 2 M8_M7_CDNS_765154963934 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X158 2 M8_M7_CDNS_765154963934 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X159 2 M8_M7_CDNS_765154963934 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X160 2 M8_M7_CDNS_765154963934 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X161 1 M8_M7_CDNS_765154963934 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X162 1 M8_M7_CDNS_765154963934 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X163 1 M8_M7_CDNS_765154963934 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X164 1 M8_M7_CDNS_765154963934 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X165 2 M8_M7_CDNS_765154963934 $T=1340 28530 0 0 $X=980 $Y=28400
X166 2 M8_M7_CDNS_765154963934 $T=1340 38870 0 0 $X=980 $Y=38740
X167 2 M8_M7_CDNS_765154963934 $T=2350 48710 0 0 $X=1990 $Y=48580
X168 2 M8_M7_CDNS_765154963934 $T=2350 58460 0 0 $X=1990 $Y=58330
X169 1 M8_M7_CDNS_765154963934 $T=6020 35670 0 0 $X=5660 $Y=35540
X170 1 M8_M7_CDNS_765154963934 $T=6020 44210 0 0 $X=5660 $Y=44080
X171 1 M8_M7_CDNS_765154963934 $T=6020 52420 0 0 $X=5660 $Y=52290
X172 1 M8_M7_CDNS_765154963934 $T=6020 62650 0 0 $X=5660 $Y=62520
X173 2 M8_M7_CDNS_765154963934 $T=7810 29790 0 0 $X=7450 $Y=29660
X174 2 M8_M7_CDNS_765154963934 $T=7810 38630 0 0 $X=7450 $Y=38500
X175 2 M8_M7_CDNS_765154963934 $T=7810 45970 0 0 $X=7450 $Y=45840
X176 2 M8_M7_CDNS_765154963934 $T=7810 54500 0 0 $X=7450 $Y=54370
X177 2 M8_M7_CDNS_765154963934 $T=23540 29510 0 0 $X=23180 $Y=29380
X178 2 M8_M7_CDNS_765154963934 $T=23540 36860 0 0 $X=23180 $Y=36730
X179 2 M8_M7_CDNS_765154963934 $T=24360 21640 0 0 $X=24000 $Y=21510
X180 2 M8_M7_CDNS_765154963934 $T=26800 45560 0 0 $X=26440 $Y=45430
X181 1 M8_M7_CDNS_765154963934 $T=28170 26920 0 0 $X=27810 $Y=26790
X182 1 M8_M7_CDNS_765154963934 $T=28170 35440 0 0 $X=27810 $Y=35310
X183 1 M8_M7_CDNS_765154963934 $T=28170 44210 0 0 $X=27810 $Y=44080
X184 1 M8_M7_CDNS_765154963934 $T=28170 53250 0 0 $X=27810 $Y=53120
X185 1 M8_M7_CDNS_765154963934 $T=28170 72500 0 0 $X=27810 $Y=72370
X186 2 M8_M7_CDNS_765154963934 $T=30470 38630 0 0 $X=30110 $Y=38500
X187 2 M8_M7_CDNS_765154963934 $T=33760 21470 0 0 $X=33400 $Y=21340
X188 2 M8_M7_CDNS_765154963934 $T=33760 29680 0 0 $X=33400 $Y=29550
X189 2 M8_M7_CDNS_765154963934 $T=34980 45870 0 0 $X=34620 $Y=45740
X190 2 M8_M7_CDNS_765154963934 $T=50880 20850 0 0 $X=50520 $Y=20720
X191 2 M8_M7_CDNS_765154963934 $T=50880 28780 0 0 $X=50520 $Y=28650
X192 2 M8_M7_CDNS_765154963934 $T=50880 36650 0 0 $X=50520 $Y=36520
X193 2 M8_M7_CDNS_765154963934 $T=51050 12420 0 0 $X=50690 $Y=12290
X194 1 M8_M7_CDNS_765154963934 $T=53300 19220 0 0 $X=52940 $Y=19090
X195 1 M8_M7_CDNS_765154963934 $T=53300 26650 0 0 $X=52940 $Y=26520
X196 1 M8_M7_CDNS_765154963934 $T=53300 35880 0 0 $X=52940 $Y=35750
X197 1 M8_M7_CDNS_765154963934 $T=55090 43020 0 0 $X=54730 $Y=42890
X198 2 M8_M7_CDNS_765154963934 $T=57390 12420 0 0 $X=57030 $Y=12290
X199 2 M8_M7_CDNS_765154963934 $T=57390 20810 0 0 $X=57030 $Y=20680
X200 2 M8_M7_CDNS_765154963934 $T=57390 29200 0 0 $X=57030 $Y=29070
X201 2 M8_M7_CDNS_765154963934 $T=57390 37590 0 0 $X=57030 $Y=37460
X202 3 M8_M7_CDNS_765154963934 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X203 2 M10_M9_CDNS_765154963935 $T=-6030 34390 0 0 $X=-6990 $Y=34110
X204 2 M10_M9_CDNS_765154963935 $T=-6030 43750 0 0 $X=-6990 $Y=43470
X205 2 M10_M9_CDNS_765154963935 $T=-6030 55310 0 0 $X=-6990 $Y=55030
X206 2 M10_M9_CDNS_765154963935 $T=-6030 65170 0 0 $X=-6990 $Y=64890
X207 1 M10_M9_CDNS_765154963935 $T=-4370 38930 0 0 $X=-5330 $Y=38650
X208 1 M10_M9_CDNS_765154963935 $T=-4370 45380 0 0 $X=-5330 $Y=45100
X209 1 M10_M9_CDNS_765154963935 $T=-4370 60080 0 0 $X=-5330 $Y=59800
X210 1 M10_M9_CDNS_765154963935 $T=-3860 70340 0 0 $X=-4820 $Y=70060
X211 2 M10_M9_CDNS_765154963935 $T=1340 28520 0 0 $X=380 $Y=28240
X212 2 M10_M9_CDNS_765154963935 $T=1340 38860 0 0 $X=380 $Y=38580
X213 2 M10_M9_CDNS_765154963935 $T=2350 48700 0 0 $X=1390 $Y=48420
X214 2 M10_M9_CDNS_765154963935 $T=2350 58450 0 0 $X=1390 $Y=58170
X215 1 M10_M9_CDNS_765154963935 $T=6020 35670 0 0 $X=5060 $Y=35390
X216 1 M10_M9_CDNS_765154963935 $T=6020 44210 0 0 $X=5060 $Y=43930
X217 1 M10_M9_CDNS_765154963935 $T=6020 52420 0 0 $X=5060 $Y=52140
X218 1 M10_M9_CDNS_765154963935 $T=6020 62650 0 0 $X=5060 $Y=62370
X219 2 M10_M9_CDNS_765154963935 $T=7810 29780 0 0 $X=6850 $Y=29500
X220 2 M10_M9_CDNS_765154963935 $T=7810 38620 0 0 $X=6850 $Y=38340
X221 2 M10_M9_CDNS_765154963935 $T=7810 45960 0 0 $X=6850 $Y=45680
X222 2 M10_M9_CDNS_765154963935 $T=7810 54490 0 0 $X=6850 $Y=54210
X223 2 M10_M9_CDNS_765154963935 $T=23540 29500 0 0 $X=22580 $Y=29220
X224 2 M10_M9_CDNS_765154963935 $T=23540 36850 0 0 $X=22580 $Y=36570
X225 2 M10_M9_CDNS_765154963935 $T=24360 21640 0 0 $X=23400 $Y=21360
X226 2 M10_M9_CDNS_765154963935 $T=26490 4150 0 0 $X=25530 $Y=3870
X227 2 M10_M9_CDNS_765154963935 $T=26730 45590 0 0 $X=25770 $Y=45310
X228 1 M10_M9_CDNS_765154963935 $T=28170 26920 0 0 $X=27210 $Y=26640
X229 1 M10_M9_CDNS_765154963935 $T=28170 35440 0 0 $X=27210 $Y=35160
X230 1 M10_M9_CDNS_765154963935 $T=28170 44210 0 0 $X=27210 $Y=43930
X231 1 M10_M9_CDNS_765154963935 $T=28170 53250 0 0 $X=27210 $Y=52970
X232 1 M10_M9_CDNS_765154963935 $T=28170 72500 0 0 $X=27210 $Y=72220
X233 2 M10_M9_CDNS_765154963935 $T=30480 38640 0 0 $X=29520 $Y=38360
X234 2 M10_M9_CDNS_765154963935 $T=33760 21510 0 0 $X=32800 $Y=21230
X235 2 M10_M9_CDNS_765154963935 $T=33760 29720 0 0 $X=32800 $Y=29440
X236 2 M10_M9_CDNS_765154963935 $T=34980 45860 0 0 $X=34020 $Y=45580
X237 2 M10_M9_CDNS_765154963935 $T=50880 20890 0 0 $X=49920 $Y=20610
X238 2 M10_M9_CDNS_765154963935 $T=50880 28820 0 0 $X=49920 $Y=28540
X239 2 M10_M9_CDNS_765154963935 $T=50880 36690 0 0 $X=49920 $Y=36410
X240 2 M10_M9_CDNS_765154963935 $T=51050 12460 0 0 $X=50090 $Y=12180
X241 1 M10_M9_CDNS_765154963935 $T=53300 19220 0 0 $X=52340 $Y=18940
X242 1 M10_M9_CDNS_765154963935 $T=53300 26650 0 0 $X=52340 $Y=26370
X243 1 M10_M9_CDNS_765154963935 $T=53300 35880 0 0 $X=52340 $Y=35600
X244 1 M10_M9_CDNS_765154963935 $T=55090 43020 0 0 $X=54130 $Y=42740
X245 2 M10_M9_CDNS_765154963935 $T=57390 12460 0 0 $X=56430 $Y=12180
X246 2 M10_M9_CDNS_765154963935 $T=57390 20850 0 0 $X=56430 $Y=20570
X247 2 M10_M9_CDNS_765154963935 $T=57390 29240 0 0 $X=56430 $Y=28960
X248 2 M10_M9_CDNS_765154963935 $T=57390 37630 0 0 $X=56430 $Y=37350
X249 3 M10_M9_CDNS_765154963935 $T=77820 -5300 0 0 $X=76860 $Y=-5580
X250 2 M9_M8_CDNS_765154963936 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X251 2 M9_M8_CDNS_765154963936 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X252 2 M9_M8_CDNS_765154963936 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X253 2 M9_M8_CDNS_765154963936 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X254 1 M9_M8_CDNS_765154963936 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X255 1 M9_M8_CDNS_765154963936 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X256 1 M9_M8_CDNS_765154963936 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X257 1 M9_M8_CDNS_765154963936 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X258 2 M9_M8_CDNS_765154963936 $T=1340 28530 0 0 $X=980 $Y=28400
X259 2 M9_M8_CDNS_765154963936 $T=1340 38870 0 0 $X=980 $Y=38740
X260 2 M9_M8_CDNS_765154963936 $T=2350 48710 0 0 $X=1990 $Y=48580
X261 2 M9_M8_CDNS_765154963936 $T=2350 58460 0 0 $X=1990 $Y=58330
X262 1 M9_M8_CDNS_765154963936 $T=6020 35670 0 0 $X=5660 $Y=35540
X263 1 M9_M8_CDNS_765154963936 $T=6020 44210 0 0 $X=5660 $Y=44080
X264 1 M9_M8_CDNS_765154963936 $T=6020 52420 0 0 $X=5660 $Y=52290
X265 1 M9_M8_CDNS_765154963936 $T=6020 62650 0 0 $X=5660 $Y=62520
X266 2 M9_M8_CDNS_765154963936 $T=7810 29790 0 0 $X=7450 $Y=29660
X267 2 M9_M8_CDNS_765154963936 $T=7810 38630 0 0 $X=7450 $Y=38500
X268 2 M9_M8_CDNS_765154963936 $T=7810 45970 0 0 $X=7450 $Y=45840
X269 2 M9_M8_CDNS_765154963936 $T=7810 54500 0 0 $X=7450 $Y=54370
X270 2 M9_M8_CDNS_765154963936 $T=23540 29510 0 0 $X=23180 $Y=29380
X271 2 M9_M8_CDNS_765154963936 $T=23540 36860 0 0 $X=23180 $Y=36730
X272 2 M9_M8_CDNS_765154963936 $T=24360 21640 0 0 $X=24000 $Y=21510
X273 2 M9_M8_CDNS_765154963936 $T=26800 45560 0 0 $X=26440 $Y=45430
X274 1 M9_M8_CDNS_765154963936 $T=28170 26920 0 0 $X=27810 $Y=26790
X275 1 M9_M8_CDNS_765154963936 $T=28170 35440 0 0 $X=27810 $Y=35310
X276 1 M9_M8_CDNS_765154963936 $T=28170 44210 0 0 $X=27810 $Y=44080
X277 1 M9_M8_CDNS_765154963936 $T=28170 53250 0 0 $X=27810 $Y=53120
X278 1 M9_M8_CDNS_765154963936 $T=28170 72500 0 0 $X=27810 $Y=72370
X279 2 M9_M8_CDNS_765154963936 $T=30470 38630 0 0 $X=30110 $Y=38500
X280 2 M9_M8_CDNS_765154963936 $T=33760 21470 0 0 $X=33400 $Y=21340
X281 2 M9_M8_CDNS_765154963936 $T=33760 29680 0 0 $X=33400 $Y=29550
X282 2 M9_M8_CDNS_765154963936 $T=34980 45870 0 0 $X=34620 $Y=45740
X283 2 M9_M8_CDNS_765154963936 $T=50880 20850 0 0 $X=50520 $Y=20720
X284 2 M9_M8_CDNS_765154963936 $T=50880 28780 0 0 $X=50520 $Y=28650
X285 2 M9_M8_CDNS_765154963936 $T=50880 36650 0 0 $X=50520 $Y=36520
X286 2 M9_M8_CDNS_765154963936 $T=51050 12420 0 0 $X=50690 $Y=12290
X287 1 M9_M8_CDNS_765154963936 $T=53300 19220 0 0 $X=52940 $Y=19090
X288 1 M9_M8_CDNS_765154963936 $T=53300 26650 0 0 $X=52940 $Y=26520
X289 1 M9_M8_CDNS_765154963936 $T=53300 35880 0 0 $X=52940 $Y=35750
X290 1 M9_M8_CDNS_765154963936 $T=55090 43020 0 0 $X=54730 $Y=42890
X291 2 M9_M8_CDNS_765154963936 $T=57390 12420 0 0 $X=57030 $Y=12290
X292 2 M9_M8_CDNS_765154963936 $T=57390 20810 0 0 $X=57030 $Y=20680
X293 2 M9_M8_CDNS_765154963936 $T=57390 29200 0 0 $X=57030 $Y=29070
X294 2 M9_M8_CDNS_765154963936 $T=57390 37590 0 0 $X=57030 $Y=37460
X295 3 M9_M8_CDNS_765154963936 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X296 2 M2_M1_CDNS_765154963937 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X297 2 M2_M1_CDNS_765154963937 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X298 2 M2_M1_CDNS_765154963937 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X299 2 M2_M1_CDNS_765154963937 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X300 1 M2_M1_CDNS_765154963937 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X301 1 M2_M1_CDNS_765154963937 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X302 1 M2_M1_CDNS_765154963937 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X303 1 M2_M1_CDNS_765154963937 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X304 2 M2_M1_CDNS_765154963937 $T=1340 28530 0 0 $X=980 $Y=28400
X305 2 M2_M1_CDNS_765154963937 $T=1340 38870 0 0 $X=980 $Y=38740
X306 2 M2_M1_CDNS_765154963937 $T=2350 48710 0 0 $X=1990 $Y=48580
X307 2 M2_M1_CDNS_765154963937 $T=2350 58460 0 0 $X=1990 $Y=58330
X308 1 M2_M1_CDNS_765154963937 $T=6020 35670 0 0 $X=5660 $Y=35540
X309 1 M2_M1_CDNS_765154963937 $T=6020 44210 0 0 $X=5660 $Y=44080
X310 1 M2_M1_CDNS_765154963937 $T=6020 52420 0 0 $X=5660 $Y=52290
X311 1 M2_M1_CDNS_765154963937 $T=6020 62650 0 0 $X=5660 $Y=62520
X312 2 M2_M1_CDNS_765154963937 $T=7810 29790 0 0 $X=7450 $Y=29660
X313 2 M2_M1_CDNS_765154963937 $T=7810 38630 0 0 $X=7450 $Y=38500
X314 2 M2_M1_CDNS_765154963937 $T=7810 45970 0 0 $X=7450 $Y=45840
X315 2 M2_M1_CDNS_765154963937 $T=7810 54500 0 0 $X=7450 $Y=54370
X316 2 M2_M1_CDNS_765154963937 $T=23540 29510 0 0 $X=23180 $Y=29380
X317 2 M2_M1_CDNS_765154963937 $T=23540 36860 0 0 $X=23180 $Y=36730
X318 2 M2_M1_CDNS_765154963937 $T=24360 21640 0 0 $X=24000 $Y=21510
X319 2 M2_M1_CDNS_765154963937 $T=26800 45560 0 0 $X=26440 $Y=45430
X320 1 M2_M1_CDNS_765154963937 $T=28170 26920 0 0 $X=27810 $Y=26790
X321 1 M2_M1_CDNS_765154963937 $T=28170 35440 0 0 $X=27810 $Y=35310
X322 1 M2_M1_CDNS_765154963937 $T=28170 44210 0 0 $X=27810 $Y=44080
X323 1 M2_M1_CDNS_765154963937 $T=28170 53250 0 0 $X=27810 $Y=53120
X324 1 M2_M1_CDNS_765154963937 $T=28170 72500 0 0 $X=27810 $Y=72370
X325 2 M2_M1_CDNS_765154963937 $T=30470 38630 0 0 $X=30110 $Y=38500
X326 2 M2_M1_CDNS_765154963937 $T=33760 21470 0 0 $X=33400 $Y=21340
X327 2 M2_M1_CDNS_765154963937 $T=33760 29680 0 0 $X=33400 $Y=29550
X328 2 M2_M1_CDNS_765154963937 $T=34980 45870 0 0 $X=34620 $Y=45740
X329 2 M2_M1_CDNS_765154963937 $T=50880 20850 0 0 $X=50520 $Y=20720
X330 2 M2_M1_CDNS_765154963937 $T=50880 28780 0 0 $X=50520 $Y=28650
X331 2 M2_M1_CDNS_765154963937 $T=50880 36650 0 0 $X=50520 $Y=36520
X332 2 M2_M1_CDNS_765154963937 $T=51050 12420 0 0 $X=50690 $Y=12290
X333 1 M2_M1_CDNS_765154963937 $T=53300 19220 0 0 $X=52940 $Y=19090
X334 1 M2_M1_CDNS_765154963937 $T=53300 26650 0 0 $X=52940 $Y=26520
X335 1 M2_M1_CDNS_765154963937 $T=53300 35880 0 0 $X=52940 $Y=35750
X336 1 M2_M1_CDNS_765154963937 $T=55090 43020 0 0 $X=54730 $Y=42890
X337 2 M2_M1_CDNS_765154963937 $T=57390 12420 0 0 $X=57030 $Y=12290
X338 2 M2_M1_CDNS_765154963937 $T=57390 20810 0 0 $X=57030 $Y=20680
X339 2 M2_M1_CDNS_765154963937 $T=57390 29200 0 0 $X=57030 $Y=29070
X340 2 M2_M1_CDNS_765154963937 $T=57390 37590 0 0 $X=57030 $Y=37460
X341 3 M2_M1_CDNS_765154963937 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X342 2 M3_M2_CDNS_765154963938 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X343 2 M3_M2_CDNS_765154963938 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X344 2 M3_M2_CDNS_765154963938 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X345 2 M3_M2_CDNS_765154963938 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X346 1 M3_M2_CDNS_765154963938 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X347 1 M3_M2_CDNS_765154963938 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X348 1 M3_M2_CDNS_765154963938 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X349 1 M3_M2_CDNS_765154963938 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X350 2 M3_M2_CDNS_765154963938 $T=1340 28530 0 0 $X=980 $Y=28400
X351 2 M3_M2_CDNS_765154963938 $T=1340 38870 0 0 $X=980 $Y=38740
X352 2 M3_M2_CDNS_765154963938 $T=2350 48710 0 0 $X=1990 $Y=48580
X353 2 M3_M2_CDNS_765154963938 $T=2350 58460 0 0 $X=1990 $Y=58330
X354 1 M3_M2_CDNS_765154963938 $T=6020 35670 0 0 $X=5660 $Y=35540
X355 1 M3_M2_CDNS_765154963938 $T=6020 44210 0 0 $X=5660 $Y=44080
X356 1 M3_M2_CDNS_765154963938 $T=6020 52420 0 0 $X=5660 $Y=52290
X357 1 M3_M2_CDNS_765154963938 $T=6020 62650 0 0 $X=5660 $Y=62520
X358 2 M3_M2_CDNS_765154963938 $T=7810 29790 0 0 $X=7450 $Y=29660
X359 2 M3_M2_CDNS_765154963938 $T=7810 38630 0 0 $X=7450 $Y=38500
X360 2 M3_M2_CDNS_765154963938 $T=7810 45970 0 0 $X=7450 $Y=45840
X361 2 M3_M2_CDNS_765154963938 $T=7810 54500 0 0 $X=7450 $Y=54370
X362 2 M3_M2_CDNS_765154963938 $T=23540 29510 0 0 $X=23180 $Y=29380
X363 2 M3_M2_CDNS_765154963938 $T=23540 36860 0 0 $X=23180 $Y=36730
X364 2 M3_M2_CDNS_765154963938 $T=24360 21640 0 0 $X=24000 $Y=21510
X365 2 M3_M2_CDNS_765154963938 $T=26800 45560 0 0 $X=26440 $Y=45430
X366 1 M3_M2_CDNS_765154963938 $T=28170 26920 0 0 $X=27810 $Y=26790
X367 1 M3_M2_CDNS_765154963938 $T=28170 35440 0 0 $X=27810 $Y=35310
X368 1 M3_M2_CDNS_765154963938 $T=28170 44210 0 0 $X=27810 $Y=44080
X369 1 M3_M2_CDNS_765154963938 $T=28170 53250 0 0 $X=27810 $Y=53120
X370 1 M3_M2_CDNS_765154963938 $T=28170 72500 0 0 $X=27810 $Y=72370
X371 2 M3_M2_CDNS_765154963938 $T=30470 38630 0 0 $X=30110 $Y=38500
X372 2 M3_M2_CDNS_765154963938 $T=33760 21470 0 0 $X=33400 $Y=21340
X373 2 M3_M2_CDNS_765154963938 $T=33760 29680 0 0 $X=33400 $Y=29550
X374 2 M3_M2_CDNS_765154963938 $T=34980 45870 0 0 $X=34620 $Y=45740
X375 2 M3_M2_CDNS_765154963938 $T=50880 20850 0 0 $X=50520 $Y=20720
X376 2 M3_M2_CDNS_765154963938 $T=50880 28780 0 0 $X=50520 $Y=28650
X377 2 M3_M2_CDNS_765154963938 $T=50880 36650 0 0 $X=50520 $Y=36520
X378 2 M3_M2_CDNS_765154963938 $T=51050 12420 0 0 $X=50690 $Y=12290
X379 1 M3_M2_CDNS_765154963938 $T=53300 19220 0 0 $X=52940 $Y=19090
X380 1 M3_M2_CDNS_765154963938 $T=53300 26650 0 0 $X=52940 $Y=26520
X381 1 M3_M2_CDNS_765154963938 $T=53300 35880 0 0 $X=52940 $Y=35750
X382 1 M3_M2_CDNS_765154963938 $T=55090 43020 0 0 $X=54730 $Y=42890
X383 2 M3_M2_CDNS_765154963938 $T=57390 12420 0 0 $X=57030 $Y=12290
X384 2 M3_M2_CDNS_765154963938 $T=57390 20810 0 0 $X=57030 $Y=20680
X385 2 M3_M2_CDNS_765154963938 $T=57390 29200 0 0 $X=57030 $Y=29070
X386 2 M3_M2_CDNS_765154963938 $T=57390 37590 0 0 $X=57030 $Y=37460
X387 3 M3_M2_CDNS_765154963938 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X388 2 M4_M3_CDNS_765154963939 $T=-6030 34400 0 0 $X=-6390 $Y=34270
X389 2 M4_M3_CDNS_765154963939 $T=-6030 43760 0 0 $X=-6390 $Y=43630
X390 2 M4_M3_CDNS_765154963939 $T=-6030 55320 0 0 $X=-6390 $Y=55190
X391 2 M4_M3_CDNS_765154963939 $T=-6030 65180 0 0 $X=-6390 $Y=65050
X392 1 M4_M3_CDNS_765154963939 $T=-4370 38930 0 0 $X=-4730 $Y=38800
X393 1 M4_M3_CDNS_765154963939 $T=-4370 45380 0 0 $X=-4730 $Y=45250
X394 1 M4_M3_CDNS_765154963939 $T=-4370 60080 0 0 $X=-4730 $Y=59950
X395 1 M4_M3_CDNS_765154963939 $T=-3860 70340 0 0 $X=-4220 $Y=70210
X396 2 M4_M3_CDNS_765154963939 $T=1340 28530 0 0 $X=980 $Y=28400
X397 2 M4_M3_CDNS_765154963939 $T=1340 38870 0 0 $X=980 $Y=38740
X398 2 M4_M3_CDNS_765154963939 $T=2350 48710 0 0 $X=1990 $Y=48580
X399 2 M4_M3_CDNS_765154963939 $T=2350 58460 0 0 $X=1990 $Y=58330
X400 1 M4_M3_CDNS_765154963939 $T=6020 35670 0 0 $X=5660 $Y=35540
X401 1 M4_M3_CDNS_765154963939 $T=6020 44210 0 0 $X=5660 $Y=44080
X402 1 M4_M3_CDNS_765154963939 $T=6020 52420 0 0 $X=5660 $Y=52290
X403 1 M4_M3_CDNS_765154963939 $T=6020 62650 0 0 $X=5660 $Y=62520
X404 2 M4_M3_CDNS_765154963939 $T=7810 29790 0 0 $X=7450 $Y=29660
X405 2 M4_M3_CDNS_765154963939 $T=7810 38630 0 0 $X=7450 $Y=38500
X406 2 M4_M3_CDNS_765154963939 $T=7810 45970 0 0 $X=7450 $Y=45840
X407 2 M4_M3_CDNS_765154963939 $T=7810 54500 0 0 $X=7450 $Y=54370
X408 2 M4_M3_CDNS_765154963939 $T=23540 29510 0 0 $X=23180 $Y=29380
X409 2 M4_M3_CDNS_765154963939 $T=23540 36860 0 0 $X=23180 $Y=36730
X410 2 M4_M3_CDNS_765154963939 $T=24360 21640 0 0 $X=24000 $Y=21510
X411 2 M4_M3_CDNS_765154963939 $T=26800 45560 0 0 $X=26440 $Y=45430
X412 1 M4_M3_CDNS_765154963939 $T=28170 26920 0 0 $X=27810 $Y=26790
X413 1 M4_M3_CDNS_765154963939 $T=28170 35440 0 0 $X=27810 $Y=35310
X414 1 M4_M3_CDNS_765154963939 $T=28170 44210 0 0 $X=27810 $Y=44080
X415 1 M4_M3_CDNS_765154963939 $T=28170 53250 0 0 $X=27810 $Y=53120
X416 1 M4_M3_CDNS_765154963939 $T=28170 72500 0 0 $X=27810 $Y=72370
X417 2 M4_M3_CDNS_765154963939 $T=30470 38630 0 0 $X=30110 $Y=38500
X418 2 M4_M3_CDNS_765154963939 $T=33760 21470 0 0 $X=33400 $Y=21340
X419 2 M4_M3_CDNS_765154963939 $T=33760 29680 0 0 $X=33400 $Y=29550
X420 2 M4_M3_CDNS_765154963939 $T=34980 45870 0 0 $X=34620 $Y=45740
X421 2 M4_M3_CDNS_765154963939 $T=50880 20850 0 0 $X=50520 $Y=20720
X422 2 M4_M3_CDNS_765154963939 $T=50880 28780 0 0 $X=50520 $Y=28650
X423 2 M4_M3_CDNS_765154963939 $T=50880 36650 0 0 $X=50520 $Y=36520
X424 2 M4_M3_CDNS_765154963939 $T=51050 12420 0 0 $X=50690 $Y=12290
X425 1 M4_M3_CDNS_765154963939 $T=53300 19220 0 0 $X=52940 $Y=19090
X426 1 M4_M3_CDNS_765154963939 $T=53300 26650 0 0 $X=52940 $Y=26520
X427 1 M4_M3_CDNS_765154963939 $T=53300 35880 0 0 $X=52940 $Y=35750
X428 1 M4_M3_CDNS_765154963939 $T=55090 43020 0 0 $X=54730 $Y=42890
X429 2 M4_M3_CDNS_765154963939 $T=57390 12420 0 0 $X=57030 $Y=12290
X430 2 M4_M3_CDNS_765154963939 $T=57390 20810 0 0 $X=57030 $Y=20680
X431 2 M4_M3_CDNS_765154963939 $T=57390 29200 0 0 $X=57030 $Y=29070
X432 2 M4_M3_CDNS_765154963939 $T=57390 37590 0 0 $X=57030 $Y=37460
X433 3 M4_M3_CDNS_765154963939 $T=77820 -5300 0 0 $X=77460 $Y=-5430
X434 4 M5_M4_CDNS_7651549639310 $T=19760 37730 0 0 $X=19680 $Y=37600
X435 5 M5_M4_CDNS_7651549639310 $T=20620 46530 0 0 $X=20540 $Y=46400
X436 4 M5_M4_CDNS_7651549639310 $T=21140 37730 0 0 $X=21060 $Y=37600
X437 6 M5_M4_CDNS_7651549639310 $T=21990 58970 0 0 $X=21910 $Y=58840
X438 5 M5_M4_CDNS_7651549639310 $T=22550 46530 0 0 $X=22470 $Y=46400
X439 6 M5_M4_CDNS_7651549639310 $T=25180 58970 0 0 $X=25100 $Y=58840
X440 7 M5_M4_CDNS_7651549639310 $T=45780 56710 0 0 $X=45700 $Y=56580
X441 7 M5_M4_CDNS_7651549639310 $T=50460 56720 0 0 $X=50380 $Y=56590
X442 6 M3_M2_CDNS_7651549639311 $T=-10530 58230 0 0 $X=-10610 $Y=57820
X443 8 M3_M2_CDNS_7651549639311 $T=-10530 68030 0 0 $X=-10610 $Y=67620
X444 4 M3_M2_CDNS_7651549639311 $T=-10230 37500 0 0 $X=-10310 $Y=37090
X445 5 M3_M2_CDNS_7651549639311 $T=-10230 46960 0 0 $X=-10310 $Y=46550
X446 9 M3_M2_CDNS_7651549639311 $T=-9230 57940 0 0 $X=-9310 $Y=57530
X447 9 M3_M2_CDNS_7651549639311 $T=-9230 67730 0 0 $X=-9310 $Y=67320
X448 9 M3_M2_CDNS_7651549639311 $T=-8930 37200 0 0 $X=-9010 $Y=36790
X449 9 M3_M2_CDNS_7651549639311 $T=-8930 46670 0 0 $X=-9010 $Y=46260
X450 4 M3_M2_CDNS_7651549639311 $T=-2010 31880 0 0 $X=-2090 $Y=31470
X451 5 M3_M2_CDNS_7651549639311 $T=-1910 42120 0 0 $X=-1990 $Y=41710
X452 6 M3_M2_CDNS_7651549639311 $T=-1910 51370 0 0 $X=-1990 $Y=50960
X453 8 M3_M2_CDNS_7651549639311 $T=-1910 61180 0 0 $X=-1990 $Y=60770
X454 10 M3_M2_CDNS_7651549639311 $T=-710 31570 0 0 $X=-790 $Y=31160
X455 10 M3_M2_CDNS_7651549639311 $T=-610 41820 0 0 $X=-690 $Y=41410
X456 10 M3_M2_CDNS_7651549639311 $T=-610 51070 0 0 $X=-690 $Y=50660
X457 10 M3_M2_CDNS_7651549639311 $T=-610 60900 0 0 $X=-690 $Y=60490
X458 4 M3_M2_CDNS_7651549639311 $T=19610 24260 0 0 $X=19530 $Y=23850
X459 5 M3_M2_CDNS_7651549639311 $T=20460 32900 0 0 $X=20380 $Y=32490
X460 11 M3_M2_CDNS_7651549639311 $T=20910 23960 0 0 $X=20830 $Y=23550
X461 6 M3_M2_CDNS_7651549639311 $T=21660 41020 0 0 $X=21580 $Y=40610
X462 11 M3_M2_CDNS_7651549639311 $T=21760 32600 0 0 $X=21680 $Y=32190
X463 11 M3_M2_CDNS_7651549639311 $T=22960 40720 0 0 $X=22880 $Y=40310
X464 8 M3_M2_CDNS_7651549639311 $T=23550 49210 0 0 $X=23470 $Y=48800
X465 11 M3_M2_CDNS_7651549639311 $T=24850 48910 0 0 $X=24770 $Y=48500
X466 4 M3_M2_CDNS_7651549639311 $T=46050 14680 0 0 $X=45970 $Y=14270
X467 5 M3_M2_CDNS_7651549639311 $T=46290 23930 0 0 $X=46210 $Y=23520
X468 6 M3_M2_CDNS_7651549639311 $T=46840 32030 0 0 $X=46760 $Y=31620
X469 12 M3_M2_CDNS_7651549639311 $T=47350 14370 0 0 $X=47270 $Y=13960
X470 12 M3_M2_CDNS_7651549639311 $T=47590 23630 0 0 $X=47510 $Y=23220
X471 12 M3_M2_CDNS_7651549639311 $T=48140 31730 0 0 $X=48060 $Y=31320
X472 8 M3_M2_CDNS_7651549639311 $T=48270 40090 0 0 $X=48190 $Y=39680
X473 12 M3_M2_CDNS_7651549639311 $T=49570 39790 0 0 $X=49490 $Y=39380
X474 6 M4_M3_CDNS_7651549639312 $T=-10530 58230 0 0 $X=-10610 $Y=57820
X475 8 M4_M3_CDNS_7651549639312 $T=-10530 68030 0 0 $X=-10610 $Y=67620
X476 4 M4_M3_CDNS_7651549639312 $T=-10230 37500 0 0 $X=-10310 $Y=37090
X477 5 M4_M3_CDNS_7651549639312 $T=-10230 46960 0 0 $X=-10310 $Y=46550
X478 4 M4_M3_CDNS_7651549639312 $T=-2010 31880 0 0 $X=-2090 $Y=31470
X479 8 M4_M3_CDNS_7651549639312 $T=-1920 61170 0 0 $X=-2000 $Y=60760
X480 5 M4_M3_CDNS_7651549639312 $T=-1910 42120 0 0 $X=-1990 $Y=41710
X481 6 M4_M3_CDNS_7651549639312 $T=-1910 51370 0 0 $X=-1990 $Y=50960
X482 4 M4_M3_CDNS_7651549639312 $T=19610 24260 0 0 $X=19530 $Y=23850
X483 5 M4_M3_CDNS_7651549639312 $T=20460 32900 0 0 $X=20380 $Y=32490
X484 6 M4_M3_CDNS_7651549639312 $T=21660 41020 0 0 $X=21580 $Y=40610
X485 8 M4_M3_CDNS_7651549639312 $T=23550 49210 0 0 $X=23470 $Y=48800
X486 4 M4_M3_CDNS_7651549639312 $T=46050 14680 0 0 $X=45970 $Y=14270
X487 5 M4_M3_CDNS_7651549639312 $T=46290 23930 0 0 $X=46210 $Y=23520
X488 6 M4_M3_CDNS_7651549639312 $T=46840 32030 0 0 $X=46760 $Y=31620
X489 8 M4_M3_CDNS_7651549639312 $T=48270 40090 0 0 $X=48190 $Y=39680
X490 6 M2_M1_CDNS_7651549639313 $T=-10530 58230 0 0 $X=-10610 $Y=57820
X491 8 M2_M1_CDNS_7651549639313 $T=-10530 68030 0 0 $X=-10610 $Y=67620
X492 4 M2_M1_CDNS_7651549639313 $T=-10230 37500 0 0 $X=-10310 $Y=37090
X493 5 M2_M1_CDNS_7651549639313 $T=-10230 46960 0 0 $X=-10310 $Y=46550
X494 9 M2_M1_CDNS_7651549639313 $T=-9230 57940 0 0 $X=-9310 $Y=57530
X495 9 M2_M1_CDNS_7651549639313 $T=-9230 67730 0 0 $X=-9310 $Y=67320
X496 9 M2_M1_CDNS_7651549639313 $T=-8930 37200 0 0 $X=-9010 $Y=36790
X497 9 M2_M1_CDNS_7651549639313 $T=-8930 46670 0 0 $X=-9010 $Y=46260
X498 4 M2_M1_CDNS_7651549639313 $T=-2010 31880 0 0 $X=-2090 $Y=31470
X499 5 M2_M1_CDNS_7651549639313 $T=-1910 42120 0 0 $X=-1990 $Y=41710
X500 6 M2_M1_CDNS_7651549639313 $T=-1910 51370 0 0 $X=-1990 $Y=50960
X501 8 M2_M1_CDNS_7651549639313 $T=-1910 61180 0 0 $X=-1990 $Y=60770
X502 10 M2_M1_CDNS_7651549639313 $T=-710 31570 0 0 $X=-790 $Y=31160
X503 10 M2_M1_CDNS_7651549639313 $T=-610 41820 0 0 $X=-690 $Y=41410
X504 10 M2_M1_CDNS_7651549639313 $T=-610 51070 0 0 $X=-690 $Y=50660
X505 10 M2_M1_CDNS_7651549639313 $T=-610 60900 0 0 $X=-690 $Y=60490
X506 4 M2_M1_CDNS_7651549639313 $T=19610 24260 0 0 $X=19530 $Y=23850
X507 5 M2_M1_CDNS_7651549639313 $T=20460 32900 0 0 $X=20380 $Y=32490
X508 11 M2_M1_CDNS_7651549639313 $T=20910 23960 0 0 $X=20830 $Y=23550
X509 6 M2_M1_CDNS_7651549639313 $T=21660 41020 0 0 $X=21580 $Y=40610
X510 11 M2_M1_CDNS_7651549639313 $T=21760 32600 0 0 $X=21680 $Y=32190
X511 11 M2_M1_CDNS_7651549639313 $T=22960 40720 0 0 $X=22880 $Y=40310
X512 8 M2_M1_CDNS_7651549639313 $T=23550 49210 0 0 $X=23470 $Y=48800
X513 11 M2_M1_CDNS_7651549639313 $T=24850 48910 0 0 $X=24770 $Y=48500
X514 4 M2_M1_CDNS_7651549639313 $T=46050 14680 0 0 $X=45970 $Y=14270
X515 5 M2_M1_CDNS_7651549639313 $T=46290 23930 0 0 $X=46210 $Y=23520
X516 6 M2_M1_CDNS_7651549639313 $T=46840 32030 0 0 $X=46760 $Y=31620
X517 12 M2_M1_CDNS_7651549639313 $T=47350 14370 0 0 $X=47270 $Y=13960
X518 12 M2_M1_CDNS_7651549639313 $T=47590 23630 0 0 $X=47510 $Y=23220
X519 12 M2_M1_CDNS_7651549639313 $T=48140 31730 0 0 $X=48060 $Y=31320
X520 8 M2_M1_CDNS_7651549639313 $T=48270 40090 0 0 $X=48190 $Y=39680
X521 12 M2_M1_CDNS_7651549639313 $T=49570 39790 0 0 $X=49490 $Y=39380
X522 13 M3_M2_CDNS_7651549639314 $T=1300 31930 0 0 $X=1220 $Y=31800
X523 14 M3_M2_CDNS_7651549639314 $T=4490 42090 0 0 $X=4410 $Y=41960
X524 15 M3_M2_CDNS_7651549639314 $T=4690 50170 0 0 $X=4610 $Y=50040
X525 16 M3_M2_CDNS_7651549639314 $T=5100 41080 0 0 $X=5020 $Y=40950
X526 17 M3_M2_CDNS_7651549639314 $T=5140 40140 0 0 $X=5060 $Y=40010
X527 18 M3_M2_CDNS_7651549639314 $T=6030 48480 0 0 $X=5950 $Y=48350
X528 19 M3_M2_CDNS_7651549639314 $T=6040 49420 0 0 $X=5960 $Y=49290
X529 20 M3_M2_CDNS_7651549639314 $T=7240 33720 0 0 $X=7160 $Y=33590
X530 21 M3_M2_CDNS_7651549639314 $T=8470 57580 0 0 $X=8390 $Y=57450
X531 22 M3_M2_CDNS_7651549639314 $T=8480 57110 0 0 $X=8400 $Y=56980
X532 23 M3_M2_CDNS_7651549639314 $T=25320 32950 0 0 $X=25240 $Y=32820
X533 24 M3_M2_CDNS_7651549639314 $T=25330 24310 0 0 $X=25250 $Y=24180
X534 25 M3_M2_CDNS_7651549639314 $T=26510 23730 0 0 $X=26430 $Y=23600
X535 26 M3_M2_CDNS_7651549639314 $T=27230 41080 0 0 $X=27150 $Y=40950
X536 27 M3_M2_CDNS_7651549639314 $T=29070 49270 0 0 $X=28990 $Y=49140
X537 28 M3_M2_CDNS_7651549639314 $T=30110 32490 0 0 $X=30030 $Y=32360
X538 29 M3_M2_CDNS_7651549639314 $T=30190 40640 0 0 $X=30110 $Y=40510
X539 30 M3_M2_CDNS_7651549639314 $T=30240 24240 0 0 $X=30160 $Y=24110
X540 31 M3_M2_CDNS_7651549639314 $T=52100 24040 0 0 $X=52020 $Y=23910
X541 32 M3_M2_CDNS_7651549639314 $T=52290 15500 0 0 $X=52210 $Y=15370
X542 33 M3_M2_CDNS_7651549639314 $T=52440 32440 0 0 $X=52360 $Y=32310
X543 34 M3_M2_CDNS_7651549639314 $T=53320 14710 0 0 $X=53240 $Y=14580
X544 35 M3_M2_CDNS_7651549639314 $T=54090 40990 0 0 $X=54010 $Y=40860
X545 36 M3_M2_CDNS_7651549639314 $T=55490 32090 0 0 $X=55410 $Y=31960
X546 37 M3_M2_CDNS_7651549639314 $T=55580 15240 0 0 $X=55500 $Y=15110
X547 38 M3_M2_CDNS_7651549639314 $T=55860 23680 0 0 $X=55780 $Y=23550
X548 22 M2_M1_CDNS_7651549639315 $T=-7220 58290 0 0 $X=-7300 $Y=58160
X549 39 M2_M1_CDNS_7651549639315 $T=-7210 68080 0 0 $X=-7290 $Y=67950
X550 17 M2_M1_CDNS_7651549639315 $T=-6920 37560 0 0 $X=-7000 $Y=37430
X551 18 M2_M1_CDNS_7651549639315 $T=-6920 47030 0 0 $X=-7000 $Y=46900
X552 13 M2_M1_CDNS_7651549639315 $T=1300 31930 0 0 $X=1220 $Y=31800
X553 19 M2_M1_CDNS_7651549639315 $T=1400 51420 0 0 $X=1320 $Y=51290
X554 21 M2_M1_CDNS_7651549639315 $T=1400 61250 0 0 $X=1320 $Y=61120
X555 16 M2_M1_CDNS_7651549639315 $T=1410 42180 0 0 $X=1330 $Y=42050
X556 24 M2_M1_CDNS_7651549639315 $T=22920 24320 0 0 $X=22840 $Y=24190
X557 23 M2_M1_CDNS_7651549639315 $T=23780 32950 0 0 $X=23700 $Y=32820
X558 26 M2_M1_CDNS_7651549639315 $T=25020 41080 0 0 $X=24940 $Y=40950
X559 27 M2_M1_CDNS_7651549639315 $T=26870 49270 0 0 $X=26790 $Y=49140
X560 32 M2_M1_CDNS_7651549639315 $T=49350 14720 0 0 $X=49270 $Y=14590
X561 31 M2_M1_CDNS_7651549639315 $T=49610 24000 0 0 $X=49530 $Y=23870
X562 33 M2_M1_CDNS_7651549639315 $T=50150 32070 0 0 $X=50070 $Y=31940
X563 35 M2_M1_CDNS_7651549639315 $T=51580 40150 0 0 $X=51500 $Y=40020
X564 4 M4_M3_CDNS_7651549639317 $T=-13540 37740 0 0 $X=-13900 $Y=37250
X565 5 M4_M3_CDNS_7651549639317 $T=-13440 46520 0 0 $X=-13800 $Y=46030
X566 6 M4_M3_CDNS_7651549639318 $T=-13520 58970 0 0 $X=-13960 $Y=58560
X567 8 M4_M3_CDNS_7651549639318 $T=-13330 68220 0 0 $X=-13770 $Y=67810
X568 40 M4_M3_CDNS_7651549639319 $T=20350 30860 0 0 $X=20270 $Y=30730
X569 41 M4_M3_CDNS_7651549639319 $T=21110 40150 0 0 $X=21030 $Y=40020
X570 42 M4_M3_CDNS_7651549639319 $T=22630 47680 0 0 $X=22550 $Y=47550
X571 7 M4_M3_CDNS_7651549639319 $T=24080 56710 0 0 $X=24000 $Y=56580
X572 40 M4_M3_CDNS_7651549639319 $T=25150 30860 0 0 $X=25070 $Y=30730
X573 41 M4_M3_CDNS_7651549639319 $T=25930 40140 0 0 $X=25850 $Y=40010
X574 42 M4_M3_CDNS_7651549639319 $T=29020 47680 0 0 $X=28940 $Y=47550
X575 43 M4_M3_CDNS_7651549639319 $T=46610 21760 0 0 $X=46530 $Y=21630
X576 44 M4_M3_CDNS_7651549639319 $T=46820 30140 0 0 $X=46740 $Y=30010
X577 45 M4_M3_CDNS_7651549639319 $T=47710 38370 0 0 $X=47630 $Y=38240
X578 46 M4_M3_CDNS_7651549639319 $T=48850 48160 0 0 $X=48770 $Y=48030
X579 43 M4_M3_CDNS_7651549639319 $T=51050 21760 0 0 $X=50970 $Y=21630
X580 44 M4_M3_CDNS_7651549639319 $T=52190 30140 0 0 $X=52110 $Y=30010
X581 45 M4_M3_CDNS_7651549639319 $T=53130 38360 0 0 $X=53050 $Y=38230
X582 46 M4_M3_CDNS_7651549639319 $T=72210 52580 0 0 $X=72130 $Y=52450
X583 7 M4_M3_CDNS_7651549639319 $T=73150 62580 0 0 $X=73070 $Y=62450
X584 6 1 9 2 22 108 52 and2 $T=-8180 57870 0 0 $X=-10850 $Y=55290
X585 8 1 9 2 39 109 53 and2 $T=-8180 67670 0 0 $X=-10850 $Y=65090
X586 4 1 9 2 17 110 54 and2 $T=-7880 37140 0 0 $X=-10550 $Y=34560
X587 5 1 9 2 18 111 55 and2 $T=-7880 46610 0 0 $X=-10550 $Y=44030
X588 4 1 10 2 13 112 56 and2 $T=340 31510 0 0 $X=-2330 $Y=28930
X589 5 1 10 2 16 113 57 and2 $T=440 41760 0 0 $X=-2230 $Y=39180
X590 6 1 10 2 19 114 58 and2 $T=440 51010 0 0 $X=-2230 $Y=48430
X591 8 1 10 2 21 115 59 and2 $T=440 60830 0 0 $X=-2230 $Y=58250
X592 4 1 11 2 24 116 60 and2 $T=21960 23900 0 0 $X=19290 $Y=21320
X593 5 1 11 2 23 117 61 and2 $T=22810 32540 0 0 $X=20140 $Y=29960
X594 6 1 11 2 26 118 62 and2 $T=24010 40660 0 0 $X=21340 $Y=38080
X595 8 1 11 2 27 119 63 and2 $T=25900 48850 0 0 $X=23230 $Y=46270
X596 4 1 12 2 32 120 64 and2 $T=48400 14310 0 0 $X=45730 $Y=11730
X597 5 1 12 2 31 121 65 and2 $T=48640 23570 0 0 $X=45970 $Y=20990
X598 6 1 12 2 33 122 66 and2 $T=49190 31670 0 0 $X=46520 $Y=29090
X599 8 1 12 2 35 123 67 and2 $T=50620 39730 0 0 $X=47950 $Y=37150
X600 16 17 14 1 2 41 20 70 69 71
+ 68 full_adder $T=4810 37240 0 0 $X=6590 $Y=38490
X601 19 18 15 1 2 42 14 74 73 75
+ 72 full_adder $T=4810 45580 0 0 $X=6590 $Y=46830
X602 23 40 28 1 2 44 30 78 77 79
+ 76 full_adder $T=29920 29020 0 0 $X=31700 $Y=30270
X603 26 41 29 1 2 45 28 82 81 83
+ 80 full_adder $T=29920 37240 0 0 $X=31700 $Y=38490
X604 24 25 30 1 2 43 34 86 85 87
+ 84 full_adder $T=30520 20800 0 0 $X=32300 $Y=22050
X605 33 44 36 1 2 47 38 90 89 91
+ 88 full_adder $T=55120 28680 0 0 $X=56900 $Y=29930
X606 31 43 38 1 2 48 37 94 93 95
+ 92 full_adder $T=55780 20220 0 0 $X=57560 $Y=21470
X607 32 34 37 1 2 49 50 98 97 99
+ 96 full_adder $T=55790 11770 0 0 $X=57570 $Y=13020
X608 20 13 2 1 40 25 100 half_adder $T=5880 29570 0 0 $X=8180 $Y=29850
X609 21 22 2 1 7 15 102 half_adder $T=6180 54010 0 0 $X=8480 $Y=54290
X610 27 42 2 1 46 29 104 half_adder $T=31290 45450 0 0 $X=33590 $Y=45730
X611 35 45 2 1 51 36 106 half_adder $T=55500 37450 0 0 $X=57800 $Y=37730
M0 52 6 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10430 $Y=58800 $dt=1
M1 53 8 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10430 $Y=68600 $dt=1
M2 54 4 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10130 $Y=38070 $dt=1
M3 55 5 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-10130 $Y=47540 $dt=1
M4 1 6 52 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-10020 $Y=58800 $dt=1
M5 1 8 53 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-10020 $Y=68600 $dt=1
M6 1 4 54 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-9720 $Y=38070 $dt=1
M7 1 5 55 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-9720 $Y=47540 $dt=1
M8 52 9 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-9130 $Y=58800 $dt=1
M9 53 9 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-9130 $Y=68600 $dt=1
M10 54 9 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-8830 $Y=38070 $dt=1
M11 55 9 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-8830 $Y=47540 $dt=1
M12 56 4 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1910 $Y=32440 $dt=1
M13 57 5 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1810 $Y=42690 $dt=1
M14 58 6 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1810 $Y=51940 $dt=1
M15 59 8 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-1810 $Y=61760 $dt=1
M16 1 4 56 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1500 $Y=32440 $dt=1
M17 1 5 57 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1400 $Y=42690 $dt=1
M18 1 6 58 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1400 $Y=51940 $dt=1
M19 1 8 59 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-1400 $Y=61760 $dt=1
M20 56 10 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-610 $Y=32440 $dt=1
M21 57 10 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-510 $Y=42690 $dt=1
M22 58 10 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-510 $Y=51940 $dt=1
M23 59 10 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-510 $Y=61760 $dt=1
M24 60 4 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=19710 $Y=24830 $dt=1
M25 1 4 60 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=20120 $Y=24830 $dt=1
M26 61 5 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=20560 $Y=33470 $dt=1
M27 1 5 61 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=20970 $Y=33470 $dt=1
M28 60 11 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=21010 $Y=24830 $dt=1
M29 62 6 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=21760 $Y=41590 $dt=1
M30 61 11 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=21860 $Y=33470 $dt=1
M31 1 6 62 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=22170 $Y=41590 $dt=1
M32 62 11 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=23060 $Y=41590 $dt=1
M33 63 8 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=23650 $Y=49780 $dt=1
M34 1 8 63 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=24060 $Y=49780 $dt=1
M35 63 11 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=24950 $Y=49780 $dt=1
M36 64 4 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=46150 $Y=15240 $dt=1
M37 65 5 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=46390 $Y=24500 $dt=1
M38 1 4 64 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=46560 $Y=15240 $dt=1
M39 1 5 65 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=46800 $Y=24500 $dt=1
M40 66 6 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=46940 $Y=32600 $dt=1
M41 1 6 66 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=47350 $Y=32600 $dt=1
M42 64 12 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=47450 $Y=15240 $dt=1
M43 65 12 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=47690 $Y=24500 $dt=1
M44 66 12 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=48240 $Y=32600 $dt=1
M45 67 8 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=48370 $Y=40660 $dt=1
M46 1 8 67 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=48780 $Y=40660 $dt=1
M47 67 12 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=49670 $Y=40660 $dt=1
.ends mult
