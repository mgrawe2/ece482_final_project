* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pipeline_mult_debug                          *
* Netlisted  : Sun Dec  7 19:43:55 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M10_M9_CDNS_765158229090                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M10_M9_CDNS_765158229090 1
** N=1 EP=1 FDC=0
.ends M10_M9_CDNS_765158229090

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_765158229091                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_765158229091 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_765158229091

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765158229092                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765158229092 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765158229092

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_765158229093                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_765158229093 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_765158229093

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M11_M10_CDNS_765158229094                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M11_M10_CDNS_765158229094 1
** N=1 EP=1 FDC=0
.ends M11_M10_CDNS_765158229094

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765158229095                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765158229095 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765158229095

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M8_M7_CDNS_765158229096                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M8_M7_CDNS_765158229096 1
** N=1 EP=1 FDC=0
.ends M8_M7_CDNS_765158229096

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765158229097                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765158229097 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765158229097

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765158229098                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765158229098 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765158229098

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M9_M8_CDNS_765158229099                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M9_M8_CDNS_765158229099 1
** N=1 EP=1 FDC=0
.ends M9_M8_CDNS_765158229099

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7651582290910                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7651582290910 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7651582290910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651582290911                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651582290911 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651582290911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651582290912                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651582290912 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651582290912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651582290913                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651582290913 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651582290913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651582290914                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651582290914 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651582290914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651582290915                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651582290915 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651582290915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651582290916                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651582290916 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651582290916

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651582290917                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651582290917 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651582290917

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651582290918                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651582290918 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651582290918

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651582290919                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651582290919 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651582290919

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651582290920                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651582290920 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651582290920

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651582290921                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651582290921 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651582290921

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_7651582290922                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_7651582290922 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_7651582290922

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651582290923                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651582290923 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651582290923

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_7651582290924                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_7651582290924 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_7651582290924

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651582290925                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651582290925 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651582290925

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158229090                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158229090 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 4 1 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=0 $Y=0 $dt=0
M1 2 4 3 5 g45n1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.60561 scb=0.000231313 scc=1.03051e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765158229090

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765158229091                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765158229091 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_765158229091

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158229092                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158229092 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_765158229092

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X0 2 M1_NWELL_CDNS_7651582290922 $T=190 2570 0 0 $X=-230 $Y=2270
X1 4 M1_PSUB_CDNS_7651582290924 $T=190 -2020 0 0 $X=-190 $Y=-2160
X2 1 M1_PO_CDNS_7651582290925 $T=-160 30 0 0 $X=-260 $Y=-330
X3 2 3 1 2 4 2 pmos1v_CDNS_765158229091 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 3 1 4 4 nmos1v_CDNS_765158229092 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=9
X0 2 M1_NWELL_CDNS_7651582290922 $T=-1350 2870 0 0 $X=-1770 $Y=2570
X1 6 M2_M1_CDNS_7651582290923 $T=-2410 -1220 0 0 $X=-2490 $Y=-1470
X2 7 M2_M1_CDNS_7651582290923 $T=-2000 1650 0 0 $X=-2080 $Y=1400
X3 6 M2_M1_CDNS_7651582290923 $T=-1590 -1220 0 0 $X=-1670 $Y=-1470
X4 6 M2_M1_CDNS_7651582290923 $T=-1110 -1220 0 0 $X=-1190 $Y=-1470
X5 7 M2_M1_CDNS_7651582290923 $T=-700 1650 0 0 $X=-780 $Y=1400
X6 6 M2_M1_CDNS_7651582290923 $T=-290 -1220 0 0 $X=-370 $Y=-1470
X7 4 M1_PSUB_CDNS_7651582290924 $T=-700 -2440 0 0 $X=-1080 $Y=-2580
X8 1 M1_PO_CDNS_7651582290925 $T=-2350 360 0 0 $X=-2450 $Y=0
X9 3 M1_PO_CDNS_7651582290925 $T=-1050 60 0 0 $X=-1150 $Y=-300
X10 6 6 7 1 4 nmos1v_CDNS_765158229090 $T=-2250 -1940 0 0 $X=-2670 $Y=-2140
X11 6 6 4 3 4 nmos1v_CDNS_765158229090 $T=-950 -1940 0 0 $X=-1370 $Y=-2140
X12 2 7 1 2 4 2 pmos1v_CDNS_765158229091 $T=-2250 930 0 0 $X=-2670 $Y=730
X13 2 7 3 2 4 2 pmos1v_CDNS_765158229091 $T=-950 930 0 0 $X=-1370 $Y=730
X14 7 2 5 4 inv $T=410 300 0 0 $X=-70 $Y=-1860
M0 2 3 7 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-540 $Y=930 $dt=1
M1 5 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=350 $Y=930 $dt=1
M2 2 7 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=760 $Y=930 $dt=1
.ends and2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651582290926                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651582290926 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651582290926

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651582290927                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651582290927 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651582290927

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651582290930                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651582290930 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651582290930

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7651582290932                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7651582290932 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7651582290932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X0 5 M2_M1_CDNS_7651582290923 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X1 5 M2_M1_CDNS_7651582290923 $T=-660 950 0 0 $X=-740 $Y=700
X2 5 M2_M1_CDNS_7651582290923 $T=160 -1560 0 0 $X=80 $Y=-1810
X3 5 M2_M1_CDNS_7651582290923 $T=160 950 0 0 $X=80 $Y=700
X4 5 M2_M1_CDNS_7651582290923 $T=1050 -1560 0 0 $X=970 $Y=-1810
X5 5 M2_M1_CDNS_7651582290923 $T=1050 950 0 0 $X=970 $Y=700
X6 5 6 1 5 3 2 pmos1v_CDNS_765158229091 $T=-500 230 0 0 $X=-920 $Y=30
X7 1 5 6 1 3 2 pmos1v_CDNS_765158229091 $T=800 230 0 0 $X=380 $Y=30
X8 5 6 4 5 3 nmos1v_CDNS_765158229092 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X9 4 5 6 4 3 nmos1v_CDNS_765158229092 $T=800 -1920 0 0 $X=380 $Y=-2120
X10 1 2 4 3 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
X11 6 M2_M1_CDNS_7651582290926 $T=-30 -450 0 0 $X=-160 $Y=-580
X12 5 M2_M1_CDNS_7651582290926 $T=1330 -190 0 0 $X=1200 $Y=-320
X13 6 M2_M1_CDNS_7651582290927 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X14 6 M2_M1_CDNS_7651582290927 $T=-250 380 0 0 $X=-380 $Y=250
X15 1 M1_PO_CDNS_7651582290930 $T=-450 10 0 0 $X=-550 $Y=-110
X16 1 M1_PO_CDNS_7651582290930 $T=-450 1890 0 0 $X=-550 $Y=1770
X17 4 M1_PO_CDNS_7651582290930 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X18 1 M1_PO_CDNS_7651582290930 $T=-40 1890 0 0 $X=-140 $Y=1770
X19 6 M1_PO_CDNS_7651582290930 $T=850 -980 0 0 $X=750 $Y=-1100
X20 4 M1_PO_CDNS_7651582290932 $T=-250 -840 0 0 $X=-470 $Y=-960
M0 5 1 6 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 5 6 1 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 1 6 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 7
** N=9 EP=7 FDC=24
X0 6 M2_M1_CDNS_7651582290914 $T=9970 3310 0 0 $X=9890 $Y=3180
X1 5 M2_M1_CDNS_7651582290914 $T=10180 2730 0 0 $X=10100 $Y=2600
X2 1 M3_M2_CDNS_7651582290915 $T=2760 3570 0 0 $X=2680 $Y=3440
X3 2 M3_M2_CDNS_7651582290915 $T=4630 3110 0 0 $X=4550 $Y=2980
X4 6 M3_M2_CDNS_7651582290915 $T=9970 3310 0 0 $X=9890 $Y=3180
X5 5 M3_M2_CDNS_7651582290915 $T=10180 2730 0 0 $X=10100 $Y=2600
X6 2 4 1 3 6 9 8 and2 $T=9010 2860 0 0 $X=6340 $Y=280
X7 1 M2_M1_CDNS_7651582290926 $T=2760 2580 0 0 $X=2630 $Y=2450
X8 1 M2_M1_CDNS_7651582290926 $T=7960 2810 0 0 $X=7830 $Y=2680
X9 5 M2_M1_CDNS_7651582290927 $T=6360 3430 0 0 $X=6230 $Y=3300
X10 1 4 3 7 5 2 xor $T=4660 3560 0 0 $X=2440 $Y=1000
M0 7 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2860 $Y=3790 $dt=1
M1 4 1 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3270 $Y=3790 $dt=1
M2 2 1 5 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4160 $Y=3790 $dt=1
M3 8 2 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6760 $Y=3790 $dt=1
M4 4 2 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7170 $Y=3790 $dt=1
M5 8 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8060 $Y=3790 $dt=1
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651582290933                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651582290933 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651582290933

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158229093                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158229093 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_765158229093

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765158229094                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765158229094 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_765158229094

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=8
X0 1 M2_M1_CDNS_7651582290914 $T=-830 -970 0 0 $X=-910 $Y=-1100
X1 2 M2_M1_CDNS_7651582290914 $T=-220 -60 0 0 $X=-300 $Y=-190
X2 2 M2_M1_CDNS_7651582290914 $T=200 730 0 0 $X=120 $Y=600
X3 1 M2_M1_CDNS_7651582290914 $T=810 -970 0 0 $X=730 $Y=-1100
X4 4 M1_NWELL_CDNS_7651582290922 $T=-10 2990 0 0 $X=-430 $Y=2690
X5 5 M1_PSUB_CDNS_7651582290924 $T=0 -1600 0 0 $X=-380 $Y=-1740
X6 3 M1_PO_CDNS_7651582290925 $T=-590 550 0 0 $X=-690 $Y=190
X7 7 M1_PO_CDNS_7651582290925 $T=570 550 0 0 $X=470 $Y=190
X8 2 M1_PO_CDNS_7651582290930 $T=-220 -60 0 0 $X=-320 $Y=-180
X9 6 M1_PO_CDNS_7651582290930 $T=-210 730 0 0 $X=-310 $Y=610
X10 6 M1_PO_CDNS_7651582290930 $T=190 -60 0 0 $X=90 $Y=-180
X11 2 M1_PO_CDNS_7651582290930 $T=200 730 0 0 $X=100 $Y=610
X12 1 8 3 5 9 2 6 1 7 nmos1v_CDNS_765158229093 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 1 10 4 3 6 11 1 2 7 5
+ 4 pmos1v_CDNS_765158229094 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder 1 2 3 4 5 6 7 8 9 10
+ 11
** N=15 EP=11 FDC=36
X0 2 M2_M1_CDNS_7651582290914 $T=5250 3070 0 0 $X=5170 $Y=2940
X1 8 M2_M1_CDNS_7651582290914 $T=9530 2380 0 0 $X=9450 $Y=2250
X2 9 M2_M1_CDNS_7651582290914 $T=9530 5090 0 0 $X=9450 $Y=4960
X3 4 M2_M1_CDNS_7651582290914 $T=10820 5970 0 0 $X=10740 $Y=5840
X4 8 M2_M1_CDNS_7651582290914 $T=11040 2940 0 0 $X=10960 $Y=2810
X5 2 M2_M1_CDNS_7651582290914 $T=11390 3320 0 0 $X=11310 $Y=3190
X6 7 M2_M1_CDNS_7651582290914 $T=12920 3510 0 0 $X=12840 $Y=3380
X7 1 M3_M2_CDNS_7651582290915 $T=2270 3860 0 0 $X=2190 $Y=3730
X8 2 M3_M2_CDNS_7651582290915 $T=5790 3080 0 0 $X=5710 $Y=2950
X9 6 M3_M2_CDNS_7651582290915 $T=9120 4760 0 0 $X=9040 $Y=4630
X10 2 M3_M2_CDNS_7651582290915 $T=11410 2940 0 0 $X=11330 $Y=2810
X11 7 M3_M2_CDNS_7651582290915 $T=12920 3510 0 0 $X=12840 $Y=3380
X12 2 M4_M3_CDNS_7651582290919 $T=6980 3080 0 0 $X=6900 $Y=2950
X13 2 M4_M3_CDNS_7651582290919 $T=10140 2970 0 0 $X=10060 $Y=2840
X14 10 4 7 5 inv $T=12350 3410 0 0 $X=11870 $Y=1250
X15 4 M2_M1_CDNS_7651582290926 $T=6470 5920 0 0 $X=6340 $Y=5790
X16 3 M2_M1_CDNS_7651582290926 $T=7620 3360 0 0 $X=7490 $Y=3230
X17 3 M2_M1_CDNS_7651582290926 $T=10320 3640 0 0 $X=10190 $Y=3510
X18 4 M2_M1_CDNS_7651582290927 $T=3420 5920 0 0 $X=3290 $Y=5790
X19 1 4 5 11 9 2 xor $T=4170 3810 0 0 $X=1950 $Y=1250
X20 9 4 5 8 6 3 xor $T=8070 3810 0 0 $X=5850 $Y=1250
X21 3 M3_M2_CDNS_7651582290933 $T=7300 3360 0 0 $X=7170 $Y=3230
X22 3 M3_M2_CDNS_7651582290933 $T=10110 3640 0 0 $X=9980 $Y=3510
X23 10 9 3 4 5 8 2 12 13 14
+ 15 fa_co_network $T=10840 2990 0 0 $X=9750 $Y=1250
M0 11 1 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=2370 $Y=4040 $dt=1
M1 4 1 11 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=2780 $Y=4040 $dt=1
M2 2 1 9 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=3670 $Y=4040 $dt=1
M3 8 9 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6270 $Y=4040 $dt=1
M4 4 9 8 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=6680 $Y=4040 $dt=1
M5 3 9 6 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7570 $Y=4040 $dt=1
M6 7 10 4 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=12290 $Y=4040 $dt=1
M7 4 10 7 4 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=12700 $Y=4040 $dt=1
.ends full_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765158229095                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765158229095 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765158229095

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158229096                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158229096 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765158229096

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765158229097                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765158229097 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_765158229097

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: c2mos                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt c2mos 1 2 3 4 5 6 7 8 11 12
*.DEVICECLIMB
** N=12 EP=10 FDC=9
X0 1 M2_M1_CDNS_7651582290914 $T=480 1970 0 90 $X=350 $Y=1890
X1 7 M2_M1_CDNS_7651582290914 $T=1070 1420 0 90 $X=940 $Y=1340
X2 1 M2_M1_CDNS_7651582290914 $T=3650 1970 0 90 $X=3520 $Y=1890
X3 7 M2_M1_CDNS_7651582290914 $T=3660 1420 0 90 $X=3530 $Y=1340
X4 8 M2_M1_CDNS_7651582290914 $T=4060 1720 0 90 $X=3930 $Y=1640
X5 8 M2_M1_CDNS_7651582290914 $T=5220 1720 0 90 $X=5090 $Y=1640
X6 1 M2_M1_CDNS_7651582290914 $T=5960 2040 0 90 $X=5830 $Y=1960
X7 7 M2_M1_CDNS_7651582290914 $T=6620 1970 0 90 $X=6490 $Y=1890
X8 1 M1_PO_CDNS_7651582290930 $T=3660 1980 0 90 $X=3540 $Y=1880
X9 7 M1_PO_CDNS_7651582290930 $T=3670 1420 0 90 $X=3550 $Y=1320
X10 8 M1_PO_CDNS_7651582290930 $T=5210 1720 0 90 $X=5090 $Y=1620
X11 7 M1_PO_CDNS_7651582290930 $T=6630 1980 0 90 $X=6510 $Y=1880
X12 1 M1_PO_CDNS_7651582290930 $T=6660 1400 0 90 $X=6540 $Y=1300
X13 1 M1_PO_CDNS_7651582290932 $T=530 1970 0 0 $X=310 $Y=1850
X14 4 M1_PO_CDNS_7651582290932 $T=2110 1720 0 0 $X=1890 $Y=1600
X15 6 M1_PO_CDNS_7651582290932 $T=8090 1590 0 0 $X=7870 $Y=1470
X16 2 7 1 3 2 pmos1v_CDNS_765158229095 $T=750 2360 0 0 $X=330 $Y=2160
X17 2 9 4 3 2 pmos1v_CDNS_765158229095 $T=2240 2360 0 0 $X=1820 $Y=2160
X18 9 8 1 3 2 pmos1v_CDNS_765158229095 $T=3740 2350 0 0 $X=3320 $Y=2150
X19 2 10 8 3 2 pmos1v_CDNS_765158229095 $T=5230 2360 0 0 $X=4810 $Y=2160
X20 10 5 7 3 2 pmos1v_CDNS_765158229095 $T=6720 2340 0 0 $X=6300 $Y=2140
X21 3 1 7 3 nmos1v_CDNS_765158229096 $T=750 650 0 0 $X=330 $Y=450
X22 3 4 11 3 nmos1v_CDNS_765158229096 $T=2240 650 0 0 $X=1820 $Y=450
X23 11 7 8 3 nmos1v_CDNS_765158229096 $T=3750 650 0 0 $X=3330 $Y=450
X24 3 8 12 3 nmos1v_CDNS_765158229096 $T=5230 650 0 0 $X=4810 $Y=450
X25 12 1 5 3 nmos1v_CDNS_765158229096 $T=6720 650 0 0 $X=6300 $Y=450
X26 5 3 6 nmos1v_CDNS_765158229097 $T=8210 170 0 0 $X=7790 $Y=-30
M0 11 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=2240 $Y=650 $dt=0
M1 8 7 11 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=3750 $Y=650 $dt=0
M2 12 8 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=5230 $Y=650 $dt=0
M3 5 1 12 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=6720 $Y=650 $dt=0
M4 7 1 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.27 scb=0.0231774 scc=0.00199917 $X=750 $Y=2360 $dt=1
M5 9 4 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=2240 $Y=2360 $dt=1
M6 8 1 9 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.7063 scb=0.016025 scc=0.00198503 $X=3740 $Y=2350 $dt=1
M7 10 8 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.8778 scb=0.0157187 scc=0.00185543 $X=5230 $Y=2360 $dt=1
M8 5 7 10 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=25.6749 scb=0.0214174 scc=0.0021813 $X=6720 $Y=2340 $dt=1
.ends c2mos

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pipeline_mult_debug                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pipeline_mult_debug 7 5 4 3 8 9 10 11 55 54
+ 53 52 59 60 61 62 63 43 2 1
** N=199 EP=20 FDC=697
X0 1 M10_M9_CDNS_765158229090 $T=-58270 -16380 0 0 $X=-59230 $Y=-16660
X1 1 M10_M9_CDNS_765158229090 $T=-58270 -7020 0 0 $X=-59230 $Y=-7300
X2 1 M10_M9_CDNS_765158229090 $T=-58270 4540 0 0 $X=-59230 $Y=4260
X3 1 M10_M9_CDNS_765158229090 $T=-58270 14400 0 0 $X=-59230 $Y=14120
X4 2 M10_M9_CDNS_765158229090 $T=-56610 -11840 0 0 $X=-57570 $Y=-12120
X5 2 M10_M9_CDNS_765158229090 $T=-56610 -5390 0 0 $X=-57570 $Y=-5670
X6 2 M10_M9_CDNS_765158229090 $T=-56610 9310 0 0 $X=-57570 $Y=9030
X7 2 M10_M9_CDNS_765158229090 $T=-56100 19570 0 0 $X=-57060 $Y=19290
X8 1 M10_M9_CDNS_765158229090 $T=-50900 -22250 0 0 $X=-51860 $Y=-22530
X9 1 M10_M9_CDNS_765158229090 $T=-50900 -11910 0 0 $X=-51860 $Y=-12190
X10 1 M10_M9_CDNS_765158229090 $T=-49890 -2070 0 0 $X=-50850 $Y=-2350
X11 1 M10_M9_CDNS_765158229090 $T=-49890 7680 0 0 $X=-50850 $Y=7400
X12 2 M10_M9_CDNS_765158229090 $T=-46220 -15100 0 0 $X=-47180 $Y=-15380
X13 2 M10_M9_CDNS_765158229090 $T=-46220 -6560 0 0 $X=-47180 $Y=-6840
X14 2 M10_M9_CDNS_765158229090 $T=-46220 1650 0 0 $X=-47180 $Y=1370
X15 2 M10_M9_CDNS_765158229090 $T=-46220 11880 0 0 $X=-47180 $Y=11600
X16 1 M10_M9_CDNS_765158229090 $T=-44430 -20990 0 0 $X=-45390 $Y=-21270
X17 1 M10_M9_CDNS_765158229090 $T=-44430 -12150 0 0 $X=-45390 $Y=-12430
X18 1 M10_M9_CDNS_765158229090 $T=-44430 -4810 0 0 $X=-45390 $Y=-5090
X19 1 M10_M9_CDNS_765158229090 $T=-44430 3720 0 0 $X=-45390 $Y=3440
X20 1 M10_M9_CDNS_765158229090 $T=-28700 -21270 0 0 $X=-29660 $Y=-21550
X21 1 M10_M9_CDNS_765158229090 $T=-28700 -13920 0 0 $X=-29660 $Y=-14200
X22 1 M10_M9_CDNS_765158229090 $T=-27880 -29130 0 0 $X=-28840 $Y=-29410
X23 1 M10_M9_CDNS_765158229090 $T=-25750 -46620 0 0 $X=-26710 $Y=-46900
X24 1 M10_M9_CDNS_765158229090 $T=-25510 -5180 0 0 $X=-26470 $Y=-5460
X25 2 M10_M9_CDNS_765158229090 $T=-24070 -23850 0 0 $X=-25030 $Y=-24130
X26 2 M10_M9_CDNS_765158229090 $T=-24070 -15330 0 0 $X=-25030 $Y=-15610
X27 2 M10_M9_CDNS_765158229090 $T=-24070 -6560 0 0 $X=-25030 $Y=-6840
X28 2 M10_M9_CDNS_765158229090 $T=-24070 2480 0 0 $X=-25030 $Y=2200
X29 2 M10_M9_CDNS_765158229090 $T=-24070 21730 0 0 $X=-25030 $Y=21450
X30 1 M10_M9_CDNS_765158229090 $T=-21760 -12130 0 0 $X=-22720 $Y=-12410
X31 1 M10_M9_CDNS_765158229090 $T=-18480 -29260 0 0 $X=-19440 $Y=-29540
X32 1 M10_M9_CDNS_765158229090 $T=-18480 -21050 0 0 $X=-19440 $Y=-21330
X33 1 M10_M9_CDNS_765158229090 $T=-17260 -4910 0 0 $X=-18220 $Y=-5190
X34 1 M10_M9_CDNS_765158229090 $T=-1360 -29880 0 0 $X=-2320 $Y=-30160
X35 1 M10_M9_CDNS_765158229090 $T=-1360 -21950 0 0 $X=-2320 $Y=-22230
X36 1 M10_M9_CDNS_765158229090 $T=-1360 -14080 0 0 $X=-2320 $Y=-14360
X37 1 M10_M9_CDNS_765158229090 $T=-1190 -38310 0 0 $X=-2150 $Y=-38590
X38 2 M10_M9_CDNS_765158229090 $T=1060 -31550 0 0 $X=100 $Y=-31830
X39 2 M10_M9_CDNS_765158229090 $T=1060 -24120 0 0 $X=100 $Y=-24400
X40 2 M10_M9_CDNS_765158229090 $T=1060 -14890 0 0 $X=100 $Y=-15170
X41 2 M10_M9_CDNS_765158229090 $T=2890 -7750 0 0 $X=1930 $Y=-8030
X42 1 M10_M9_CDNS_765158229090 $T=7430 -37060 0 0 $X=6470 $Y=-37340
X43 1 M10_M9_CDNS_765158229090 $T=9050 -29210 0 0 $X=8090 $Y=-29490
X44 1 M10_M9_CDNS_765158229090 $T=9050 -19860 0 0 $X=8090 $Y=-20140
X45 1 M10_M9_CDNS_765158229090 $T=9050 -13080 0 0 $X=8090 $Y=-13360
X46 2 M10_M9_CDNS_765158229090 $T=23880 13850 0 0 $X=22920 $Y=13570
X47 2 M10_M9_CDNS_765158229090 $T=24550 3710 0 0 $X=23590 $Y=3430
X48 2 M10_M9_CDNS_765158229090 $T=26060 -34250 0 0 $X=25100 $Y=-34530
X49 2 M10_M9_CDNS_765158229090 $T=26060 -26210 0 0 $X=25100 $Y=-26490
X50 2 M10_M9_CDNS_765158229090 $T=26060 -19020 0 0 $X=25100 $Y=-19300
X51 2 M10_M9_CDNS_765158229090 $T=26060 -9950 0 0 $X=25100 $Y=-10230
X52 2 M10_M9_CDNS_765158229090 $T=29710 19070 0 0 $X=28750 $Y=18790
X53 1 M10_M9_CDNS_765158229090 $T=30630 -38310 0 0 $X=29670 $Y=-38590
X54 1 M10_M9_CDNS_765158229090 $T=30630 -29920 0 0 $X=29670 $Y=-30200
X55 1 M10_M9_CDNS_765158229090 $T=30630 -21530 0 0 $X=29670 $Y=-21810
X56 1 M10_M9_CDNS_765158229090 $T=30630 -13140 0 0 $X=29670 $Y=-13420
X57 1 M10_M9_CDNS_765158229090 $T=30630 -2160 0 0 $X=29670 $Y=-2440
X58 1 M10_M9_CDNS_765158229090 $T=30630 7720 0 0 $X=29670 $Y=7440
X59 1 M10_M9_CDNS_765158229090 $T=30630 13170 0 0 $X=29670 $Y=12890
X60 1 M6_M5_CDNS_765158229091 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X61 1 M6_M5_CDNS_765158229091 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X62 1 M6_M5_CDNS_765158229091 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X63 1 M6_M5_CDNS_765158229091 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X64 2 M6_M5_CDNS_765158229091 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X65 2 M6_M5_CDNS_765158229091 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X66 2 M6_M5_CDNS_765158229091 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X67 2 M6_M5_CDNS_765158229091 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X68 1 M6_M5_CDNS_765158229091 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X69 1 M6_M5_CDNS_765158229091 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X70 1 M6_M5_CDNS_765158229091 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X71 1 M6_M5_CDNS_765158229091 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X72 2 M6_M5_CDNS_765158229091 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X73 2 M6_M5_CDNS_765158229091 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X74 2 M6_M5_CDNS_765158229091 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X75 2 M6_M5_CDNS_765158229091 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X76 1 M6_M5_CDNS_765158229091 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X77 1 M6_M5_CDNS_765158229091 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X78 1 M6_M5_CDNS_765158229091 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X79 1 M6_M5_CDNS_765158229091 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X80 1 M6_M5_CDNS_765158229091 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X81 1 M6_M5_CDNS_765158229091 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X82 1 M6_M5_CDNS_765158229091 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X83 1 M6_M5_CDNS_765158229091 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X84 2 M6_M5_CDNS_765158229091 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X85 2 M6_M5_CDNS_765158229091 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X86 2 M6_M5_CDNS_765158229091 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X87 2 M6_M5_CDNS_765158229091 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X88 2 M6_M5_CDNS_765158229091 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X89 1 M6_M5_CDNS_765158229091 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X90 1 M6_M5_CDNS_765158229091 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X91 1 M6_M5_CDNS_765158229091 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X92 1 M6_M5_CDNS_765158229091 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X93 1 M6_M5_CDNS_765158229091 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X94 1 M6_M5_CDNS_765158229091 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X95 1 M6_M5_CDNS_765158229091 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X96 1 M6_M5_CDNS_765158229091 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X97 2 M6_M5_CDNS_765158229091 $T=1060 -31550 0 0 $X=700 $Y=-31680
X98 2 M6_M5_CDNS_765158229091 $T=1060 -24120 0 0 $X=700 $Y=-24250
X99 2 M6_M5_CDNS_765158229091 $T=1060 -14890 0 0 $X=700 $Y=-15020
X100 2 M6_M5_CDNS_765158229091 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X101 1 M6_M5_CDNS_765158229091 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X102 1 M6_M5_CDNS_765158229091 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X103 1 M6_M5_CDNS_765158229091 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X104 1 M6_M5_CDNS_765158229091 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X105 2 M6_M5_CDNS_765158229091 $T=23880 13850 0 0 $X=23520 $Y=13720
X106 2 M6_M5_CDNS_765158229091 $T=24550 3710 0 0 $X=24190 $Y=3580
X107 2 M6_M5_CDNS_765158229091 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X108 2 M6_M5_CDNS_765158229091 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X109 2 M6_M5_CDNS_765158229091 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X110 2 M6_M5_CDNS_765158229091 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X111 2 M6_M5_CDNS_765158229091 $T=29710 19070 0 0 $X=29350 $Y=18940
X112 1 M6_M5_CDNS_765158229091 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X113 1 M6_M5_CDNS_765158229091 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X114 1 M6_M5_CDNS_765158229091 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X115 1 M6_M5_CDNS_765158229091 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X116 1 M6_M5_CDNS_765158229091 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X117 1 M6_M5_CDNS_765158229091 $T=30630 7680 0 0 $X=30270 $Y=7550
X118 1 M6_M5_CDNS_765158229091 $T=30630 13130 0 0 $X=30270 $Y=13000
X119 1 M5_M4_CDNS_765158229092 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X120 1 M5_M4_CDNS_765158229092 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X121 1 M5_M4_CDNS_765158229092 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X122 1 M5_M4_CDNS_765158229092 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X123 2 M5_M4_CDNS_765158229092 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X124 2 M5_M4_CDNS_765158229092 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X125 2 M5_M4_CDNS_765158229092 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X126 2 M5_M4_CDNS_765158229092 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X127 1 M5_M4_CDNS_765158229092 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X128 1 M5_M4_CDNS_765158229092 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X129 1 M5_M4_CDNS_765158229092 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X130 1 M5_M4_CDNS_765158229092 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X131 2 M5_M4_CDNS_765158229092 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X132 2 M5_M4_CDNS_765158229092 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X133 2 M5_M4_CDNS_765158229092 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X134 2 M5_M4_CDNS_765158229092 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X135 1 M5_M4_CDNS_765158229092 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X136 1 M5_M4_CDNS_765158229092 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X137 1 M5_M4_CDNS_765158229092 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X138 1 M5_M4_CDNS_765158229092 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X139 1 M5_M4_CDNS_765158229092 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X140 1 M5_M4_CDNS_765158229092 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X141 1 M5_M4_CDNS_765158229092 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X142 1 M5_M4_CDNS_765158229092 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X143 2 M5_M4_CDNS_765158229092 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X144 2 M5_M4_CDNS_765158229092 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X145 2 M5_M4_CDNS_765158229092 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X146 2 M5_M4_CDNS_765158229092 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X147 2 M5_M4_CDNS_765158229092 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X148 1 M5_M4_CDNS_765158229092 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X149 1 M5_M4_CDNS_765158229092 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X150 1 M5_M4_CDNS_765158229092 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X151 1 M5_M4_CDNS_765158229092 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X152 1 M5_M4_CDNS_765158229092 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X153 1 M5_M4_CDNS_765158229092 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X154 1 M5_M4_CDNS_765158229092 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X155 1 M5_M4_CDNS_765158229092 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X156 2 M5_M4_CDNS_765158229092 $T=1060 -31550 0 0 $X=700 $Y=-31680
X157 2 M5_M4_CDNS_765158229092 $T=1060 -24120 0 0 $X=700 $Y=-24250
X158 2 M5_M4_CDNS_765158229092 $T=1060 -14890 0 0 $X=700 $Y=-15020
X159 2 M5_M4_CDNS_765158229092 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X160 1 M5_M4_CDNS_765158229092 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X161 1 M5_M4_CDNS_765158229092 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X162 1 M5_M4_CDNS_765158229092 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X163 1 M5_M4_CDNS_765158229092 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X164 2 M5_M4_CDNS_765158229092 $T=23880 13850 0 0 $X=23520 $Y=13720
X165 2 M5_M4_CDNS_765158229092 $T=24550 3710 0 0 $X=24190 $Y=3580
X166 2 M5_M4_CDNS_765158229092 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X167 2 M5_M4_CDNS_765158229092 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X168 2 M5_M4_CDNS_765158229092 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X169 2 M5_M4_CDNS_765158229092 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X170 2 M5_M4_CDNS_765158229092 $T=29710 19070 0 0 $X=29350 $Y=18940
X171 1 M5_M4_CDNS_765158229092 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X172 1 M5_M4_CDNS_765158229092 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X173 1 M5_M4_CDNS_765158229092 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X174 1 M5_M4_CDNS_765158229092 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X175 1 M5_M4_CDNS_765158229092 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X176 1 M5_M4_CDNS_765158229092 $T=30630 7680 0 0 $X=30270 $Y=7550
X177 1 M5_M4_CDNS_765158229092 $T=30630 13130 0 0 $X=30270 $Y=13000
X178 1 M7_M6_CDNS_765158229093 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X179 1 M7_M6_CDNS_765158229093 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X180 1 M7_M6_CDNS_765158229093 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X181 1 M7_M6_CDNS_765158229093 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X182 2 M7_M6_CDNS_765158229093 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X183 2 M7_M6_CDNS_765158229093 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X184 2 M7_M6_CDNS_765158229093 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X185 2 M7_M6_CDNS_765158229093 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X186 1 M7_M6_CDNS_765158229093 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X187 1 M7_M6_CDNS_765158229093 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X188 1 M7_M6_CDNS_765158229093 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X189 1 M7_M6_CDNS_765158229093 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X190 2 M7_M6_CDNS_765158229093 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X191 2 M7_M6_CDNS_765158229093 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X192 2 M7_M6_CDNS_765158229093 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X193 2 M7_M6_CDNS_765158229093 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X194 1 M7_M6_CDNS_765158229093 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X195 1 M7_M6_CDNS_765158229093 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X196 1 M7_M6_CDNS_765158229093 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X197 1 M7_M6_CDNS_765158229093 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X198 1 M7_M6_CDNS_765158229093 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X199 1 M7_M6_CDNS_765158229093 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X200 1 M7_M6_CDNS_765158229093 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X201 1 M7_M6_CDNS_765158229093 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X202 2 M7_M6_CDNS_765158229093 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X203 2 M7_M6_CDNS_765158229093 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X204 2 M7_M6_CDNS_765158229093 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X205 2 M7_M6_CDNS_765158229093 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X206 2 M7_M6_CDNS_765158229093 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X207 1 M7_M6_CDNS_765158229093 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X208 1 M7_M6_CDNS_765158229093 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X209 1 M7_M6_CDNS_765158229093 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X210 1 M7_M6_CDNS_765158229093 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X211 1 M7_M6_CDNS_765158229093 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X212 1 M7_M6_CDNS_765158229093 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X213 1 M7_M6_CDNS_765158229093 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X214 1 M7_M6_CDNS_765158229093 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X215 2 M7_M6_CDNS_765158229093 $T=1060 -31550 0 0 $X=700 $Y=-31680
X216 2 M7_M6_CDNS_765158229093 $T=1060 -24120 0 0 $X=700 $Y=-24250
X217 2 M7_M6_CDNS_765158229093 $T=1060 -14890 0 0 $X=700 $Y=-15020
X218 2 M7_M6_CDNS_765158229093 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X219 1 M7_M6_CDNS_765158229093 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X220 1 M7_M6_CDNS_765158229093 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X221 1 M7_M6_CDNS_765158229093 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X222 1 M7_M6_CDNS_765158229093 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X223 2 M7_M6_CDNS_765158229093 $T=23880 13850 0 0 $X=23520 $Y=13720
X224 2 M7_M6_CDNS_765158229093 $T=24550 3710 0 0 $X=24190 $Y=3580
X225 2 M7_M6_CDNS_765158229093 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X226 2 M7_M6_CDNS_765158229093 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X227 2 M7_M6_CDNS_765158229093 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X228 2 M7_M6_CDNS_765158229093 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X229 2 M7_M6_CDNS_765158229093 $T=29710 19070 0 0 $X=29350 $Y=18940
X230 1 M7_M6_CDNS_765158229093 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X231 1 M7_M6_CDNS_765158229093 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X232 1 M7_M6_CDNS_765158229093 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X233 1 M7_M6_CDNS_765158229093 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X234 1 M7_M6_CDNS_765158229093 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X235 1 M7_M6_CDNS_765158229093 $T=30630 7680 0 0 $X=30270 $Y=7550
X236 1 M7_M6_CDNS_765158229093 $T=30630 13130 0 0 $X=30270 $Y=13000
X237 2 M11_M10_CDNS_765158229094 $T=-56610 -11840 0 0 $X=-57570 $Y=-12120
X238 2 M11_M10_CDNS_765158229094 $T=-56610 -5390 0 0 $X=-57570 $Y=-5670
X239 2 M11_M10_CDNS_765158229094 $T=-56610 9310 0 0 $X=-57570 $Y=9030
X240 2 M11_M10_CDNS_765158229094 $T=-56100 19570 0 0 $X=-57060 $Y=19290
X241 2 M11_M10_CDNS_765158229094 $T=-46220 -15100 0 0 $X=-47180 $Y=-15380
X242 2 M11_M10_CDNS_765158229094 $T=-46220 -6560 0 0 $X=-47180 $Y=-6840
X243 2 M11_M10_CDNS_765158229094 $T=-46220 1650 0 0 $X=-47180 $Y=1370
X244 2 M11_M10_CDNS_765158229094 $T=-46220 11880 0 0 $X=-47180 $Y=11600
X245 1 M11_M10_CDNS_765158229094 $T=-25750 -46620 0 0 $X=-26710 $Y=-46900
X246 2 M11_M10_CDNS_765158229094 $T=-24070 -23850 0 0 $X=-25030 $Y=-24130
X247 2 M11_M10_CDNS_765158229094 $T=-24070 -15330 0 0 $X=-25030 $Y=-15610
X248 2 M11_M10_CDNS_765158229094 $T=-24070 -6560 0 0 $X=-25030 $Y=-6840
X249 2 M11_M10_CDNS_765158229094 $T=-24070 2480 0 0 $X=-25030 $Y=2200
X250 2 M11_M10_CDNS_765158229094 $T=-24070 21730 0 0 $X=-25030 $Y=21450
X251 2 M11_M10_CDNS_765158229094 $T=1060 -31550 0 0 $X=100 $Y=-31830
X252 2 M11_M10_CDNS_765158229094 $T=1060 -24120 0 0 $X=100 $Y=-24400
X253 2 M11_M10_CDNS_765158229094 $T=1060 -14890 0 0 $X=100 $Y=-15170
X254 2 M11_M10_CDNS_765158229094 $T=2890 -7750 0 0 $X=1930 $Y=-8030
X255 2 M11_M10_CDNS_765158229094 $T=23880 13850 0 0 $X=22920 $Y=13570
X256 2 M11_M10_CDNS_765158229094 $T=24550 3710 0 0 $X=23590 $Y=3430
X257 2 M11_M10_CDNS_765158229094 $T=26060 -34250 0 0 $X=25100 $Y=-34530
X258 2 M11_M10_CDNS_765158229094 $T=26060 -26210 0 0 $X=25100 $Y=-26490
X259 2 M11_M10_CDNS_765158229094 $T=26060 -19020 0 0 $X=25100 $Y=-19300
X260 2 M11_M10_CDNS_765158229094 $T=26060 -9950 0 0 $X=25100 $Y=-10230
X261 2 M11_M10_CDNS_765158229094 $T=29710 19070 0 0 $X=28750 $Y=18790
X262 1 M4_M3_CDNS_765158229095 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X263 1 M4_M3_CDNS_765158229095 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X264 1 M4_M3_CDNS_765158229095 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X265 1 M4_M3_CDNS_765158229095 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X266 2 M4_M3_CDNS_765158229095 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X267 2 M4_M3_CDNS_765158229095 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X268 2 M4_M3_CDNS_765158229095 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X269 2 M4_M3_CDNS_765158229095 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X270 1 M4_M3_CDNS_765158229095 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X271 1 M4_M3_CDNS_765158229095 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X272 1 M4_M3_CDNS_765158229095 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X273 1 M4_M3_CDNS_765158229095 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X274 2 M4_M3_CDNS_765158229095 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X275 2 M4_M3_CDNS_765158229095 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X276 2 M4_M3_CDNS_765158229095 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X277 2 M4_M3_CDNS_765158229095 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X278 1 M4_M3_CDNS_765158229095 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X279 1 M4_M3_CDNS_765158229095 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X280 1 M4_M3_CDNS_765158229095 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X281 1 M4_M3_CDNS_765158229095 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X282 1 M4_M3_CDNS_765158229095 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X283 1 M4_M3_CDNS_765158229095 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X284 1 M4_M3_CDNS_765158229095 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X285 1 M4_M3_CDNS_765158229095 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X286 2 M4_M3_CDNS_765158229095 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X287 2 M4_M3_CDNS_765158229095 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X288 2 M4_M3_CDNS_765158229095 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X289 2 M4_M3_CDNS_765158229095 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X290 2 M4_M3_CDNS_765158229095 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X291 1 M4_M3_CDNS_765158229095 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X292 1 M4_M3_CDNS_765158229095 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X293 1 M4_M3_CDNS_765158229095 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X294 1 M4_M3_CDNS_765158229095 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X295 1 M4_M3_CDNS_765158229095 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X296 1 M4_M3_CDNS_765158229095 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X297 1 M4_M3_CDNS_765158229095 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X298 1 M4_M3_CDNS_765158229095 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X299 2 M4_M3_CDNS_765158229095 $T=1060 -31550 0 0 $X=700 $Y=-31680
X300 2 M4_M3_CDNS_765158229095 $T=1060 -24120 0 0 $X=700 $Y=-24250
X301 2 M4_M3_CDNS_765158229095 $T=1060 -14890 0 0 $X=700 $Y=-15020
X302 2 M4_M3_CDNS_765158229095 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X303 1 M4_M3_CDNS_765158229095 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X304 1 M4_M3_CDNS_765158229095 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X305 1 M4_M3_CDNS_765158229095 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X306 1 M4_M3_CDNS_765158229095 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X307 2 M4_M3_CDNS_765158229095 $T=23880 13850 0 0 $X=23520 $Y=13720
X308 2 M4_M3_CDNS_765158229095 $T=24550 3710 0 0 $X=24190 $Y=3580
X309 2 M4_M3_CDNS_765158229095 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X310 2 M4_M3_CDNS_765158229095 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X311 2 M4_M3_CDNS_765158229095 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X312 2 M4_M3_CDNS_765158229095 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X313 2 M4_M3_CDNS_765158229095 $T=29710 19070 0 0 $X=29350 $Y=18940
X314 1 M4_M3_CDNS_765158229095 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X315 1 M4_M3_CDNS_765158229095 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X316 1 M4_M3_CDNS_765158229095 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X317 1 M4_M3_CDNS_765158229095 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X318 1 M4_M3_CDNS_765158229095 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X319 1 M4_M3_CDNS_765158229095 $T=30630 7680 0 0 $X=30270 $Y=7550
X320 1 M4_M3_CDNS_765158229095 $T=30630 13130 0 0 $X=30270 $Y=13000
X321 1 M8_M7_CDNS_765158229096 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X322 1 M8_M7_CDNS_765158229096 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X323 1 M8_M7_CDNS_765158229096 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X324 1 M8_M7_CDNS_765158229096 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X325 2 M8_M7_CDNS_765158229096 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X326 2 M8_M7_CDNS_765158229096 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X327 2 M8_M7_CDNS_765158229096 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X328 2 M8_M7_CDNS_765158229096 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X329 1 M8_M7_CDNS_765158229096 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X330 1 M8_M7_CDNS_765158229096 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X331 1 M8_M7_CDNS_765158229096 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X332 1 M8_M7_CDNS_765158229096 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X333 2 M8_M7_CDNS_765158229096 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X334 2 M8_M7_CDNS_765158229096 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X335 2 M8_M7_CDNS_765158229096 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X336 2 M8_M7_CDNS_765158229096 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X337 1 M8_M7_CDNS_765158229096 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X338 1 M8_M7_CDNS_765158229096 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X339 1 M8_M7_CDNS_765158229096 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X340 1 M8_M7_CDNS_765158229096 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X341 1 M8_M7_CDNS_765158229096 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X342 1 M8_M7_CDNS_765158229096 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X343 1 M8_M7_CDNS_765158229096 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X344 1 M8_M7_CDNS_765158229096 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X345 2 M8_M7_CDNS_765158229096 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X346 2 M8_M7_CDNS_765158229096 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X347 2 M8_M7_CDNS_765158229096 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X348 2 M8_M7_CDNS_765158229096 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X349 2 M8_M7_CDNS_765158229096 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X350 1 M8_M7_CDNS_765158229096 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X351 1 M8_M7_CDNS_765158229096 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X352 1 M8_M7_CDNS_765158229096 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X353 1 M8_M7_CDNS_765158229096 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X354 1 M8_M7_CDNS_765158229096 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X355 1 M8_M7_CDNS_765158229096 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X356 1 M8_M7_CDNS_765158229096 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X357 1 M8_M7_CDNS_765158229096 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X358 2 M8_M7_CDNS_765158229096 $T=1060 -31550 0 0 $X=700 $Y=-31680
X359 2 M8_M7_CDNS_765158229096 $T=1060 -24120 0 0 $X=700 $Y=-24250
X360 2 M8_M7_CDNS_765158229096 $T=1060 -14890 0 0 $X=700 $Y=-15020
X361 2 M8_M7_CDNS_765158229096 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X362 1 M8_M7_CDNS_765158229096 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X363 1 M8_M7_CDNS_765158229096 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X364 1 M8_M7_CDNS_765158229096 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X365 1 M8_M7_CDNS_765158229096 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X366 2 M8_M7_CDNS_765158229096 $T=23880 13850 0 0 $X=23520 $Y=13720
X367 2 M8_M7_CDNS_765158229096 $T=24550 3710 0 0 $X=24190 $Y=3580
X368 2 M8_M7_CDNS_765158229096 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X369 2 M8_M7_CDNS_765158229096 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X370 2 M8_M7_CDNS_765158229096 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X371 2 M8_M7_CDNS_765158229096 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X372 2 M8_M7_CDNS_765158229096 $T=29710 19070 0 0 $X=29350 $Y=18940
X373 1 M8_M7_CDNS_765158229096 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X374 1 M8_M7_CDNS_765158229096 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X375 1 M8_M7_CDNS_765158229096 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X376 1 M8_M7_CDNS_765158229096 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X377 1 M8_M7_CDNS_765158229096 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X378 1 M8_M7_CDNS_765158229096 $T=30630 7680 0 0 $X=30270 $Y=7550
X379 1 M8_M7_CDNS_765158229096 $T=30630 13130 0 0 $X=30270 $Y=13000
X380 1 M3_M2_CDNS_765158229097 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X381 1 M3_M2_CDNS_765158229097 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X382 1 M3_M2_CDNS_765158229097 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X383 1 M3_M2_CDNS_765158229097 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X384 2 M3_M2_CDNS_765158229097 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X385 2 M3_M2_CDNS_765158229097 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X386 2 M3_M2_CDNS_765158229097 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X387 2 M3_M2_CDNS_765158229097 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X388 1 M3_M2_CDNS_765158229097 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X389 1 M3_M2_CDNS_765158229097 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X390 1 M3_M2_CDNS_765158229097 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X391 1 M3_M2_CDNS_765158229097 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X392 2 M3_M2_CDNS_765158229097 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X393 2 M3_M2_CDNS_765158229097 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X394 2 M3_M2_CDNS_765158229097 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X395 2 M3_M2_CDNS_765158229097 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X396 1 M3_M2_CDNS_765158229097 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X397 1 M3_M2_CDNS_765158229097 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X398 1 M3_M2_CDNS_765158229097 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X399 1 M3_M2_CDNS_765158229097 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X400 1 M3_M2_CDNS_765158229097 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X401 1 M3_M2_CDNS_765158229097 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X402 1 M3_M2_CDNS_765158229097 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X403 1 M3_M2_CDNS_765158229097 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X404 2 M3_M2_CDNS_765158229097 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X405 2 M3_M2_CDNS_765158229097 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X406 2 M3_M2_CDNS_765158229097 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X407 2 M3_M2_CDNS_765158229097 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X408 2 M3_M2_CDNS_765158229097 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X409 1 M3_M2_CDNS_765158229097 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X410 1 M3_M2_CDNS_765158229097 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X411 1 M3_M2_CDNS_765158229097 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X412 1 M3_M2_CDNS_765158229097 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X413 1 M3_M2_CDNS_765158229097 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X414 1 M3_M2_CDNS_765158229097 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X415 1 M3_M2_CDNS_765158229097 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X416 1 M3_M2_CDNS_765158229097 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X417 2 M3_M2_CDNS_765158229097 $T=1060 -31550 0 0 $X=700 $Y=-31680
X418 2 M3_M2_CDNS_765158229097 $T=1060 -24120 0 0 $X=700 $Y=-24250
X419 2 M3_M2_CDNS_765158229097 $T=1060 -14890 0 0 $X=700 $Y=-15020
X420 2 M3_M2_CDNS_765158229097 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X421 1 M3_M2_CDNS_765158229097 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X422 1 M3_M2_CDNS_765158229097 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X423 1 M3_M2_CDNS_765158229097 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X424 1 M3_M2_CDNS_765158229097 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X425 2 M3_M2_CDNS_765158229097 $T=23880 13850 0 0 $X=23520 $Y=13720
X426 2 M3_M2_CDNS_765158229097 $T=24550 3710 0 0 $X=24190 $Y=3580
X427 2 M3_M2_CDNS_765158229097 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X428 2 M3_M2_CDNS_765158229097 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X429 2 M3_M2_CDNS_765158229097 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X430 2 M3_M2_CDNS_765158229097 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X431 2 M3_M2_CDNS_765158229097 $T=29710 19070 0 0 $X=29350 $Y=18940
X432 1 M3_M2_CDNS_765158229097 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X433 1 M3_M2_CDNS_765158229097 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X434 1 M3_M2_CDNS_765158229097 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X435 1 M3_M2_CDNS_765158229097 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X436 1 M3_M2_CDNS_765158229097 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X437 1 M3_M2_CDNS_765158229097 $T=30630 7680 0 0 $X=30270 $Y=7550
X438 1 M3_M2_CDNS_765158229097 $T=30630 13130 0 0 $X=30270 $Y=13000
X439 1 M2_M1_CDNS_765158229098 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X440 1 M2_M1_CDNS_765158229098 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X441 1 M2_M1_CDNS_765158229098 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X442 1 M2_M1_CDNS_765158229098 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X443 2 M2_M1_CDNS_765158229098 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X444 2 M2_M1_CDNS_765158229098 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X445 2 M2_M1_CDNS_765158229098 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X446 2 M2_M1_CDNS_765158229098 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X447 1 M2_M1_CDNS_765158229098 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X448 1 M2_M1_CDNS_765158229098 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X449 1 M2_M1_CDNS_765158229098 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X450 1 M2_M1_CDNS_765158229098 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X451 2 M2_M1_CDNS_765158229098 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X452 2 M2_M1_CDNS_765158229098 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X453 2 M2_M1_CDNS_765158229098 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X454 2 M2_M1_CDNS_765158229098 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X455 1 M2_M1_CDNS_765158229098 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X456 1 M2_M1_CDNS_765158229098 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X457 1 M2_M1_CDNS_765158229098 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X458 1 M2_M1_CDNS_765158229098 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X459 1 M2_M1_CDNS_765158229098 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X460 1 M2_M1_CDNS_765158229098 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X461 1 M2_M1_CDNS_765158229098 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X462 1 M2_M1_CDNS_765158229098 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X463 2 M2_M1_CDNS_765158229098 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X464 2 M2_M1_CDNS_765158229098 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X465 2 M2_M1_CDNS_765158229098 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X466 2 M2_M1_CDNS_765158229098 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X467 2 M2_M1_CDNS_765158229098 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X468 1 M2_M1_CDNS_765158229098 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X469 1 M2_M1_CDNS_765158229098 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X470 1 M2_M1_CDNS_765158229098 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X471 1 M2_M1_CDNS_765158229098 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X472 1 M2_M1_CDNS_765158229098 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X473 1 M2_M1_CDNS_765158229098 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X474 1 M2_M1_CDNS_765158229098 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X475 1 M2_M1_CDNS_765158229098 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X476 2 M2_M1_CDNS_765158229098 $T=1060 -31550 0 0 $X=700 $Y=-31680
X477 2 M2_M1_CDNS_765158229098 $T=1060 -24120 0 0 $X=700 $Y=-24250
X478 2 M2_M1_CDNS_765158229098 $T=1060 -14890 0 0 $X=700 $Y=-15020
X479 2 M2_M1_CDNS_765158229098 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X480 1 M2_M1_CDNS_765158229098 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X481 1 M2_M1_CDNS_765158229098 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X482 1 M2_M1_CDNS_765158229098 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X483 1 M2_M1_CDNS_765158229098 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X484 2 M2_M1_CDNS_765158229098 $T=23880 13850 0 0 $X=23520 $Y=13720
X485 2 M2_M1_CDNS_765158229098 $T=24550 3710 0 0 $X=24190 $Y=3580
X486 2 M2_M1_CDNS_765158229098 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X487 2 M2_M1_CDNS_765158229098 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X488 2 M2_M1_CDNS_765158229098 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X489 2 M2_M1_CDNS_765158229098 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X490 2 M2_M1_CDNS_765158229098 $T=29710 19070 0 0 $X=29350 $Y=18940
X491 1 M2_M1_CDNS_765158229098 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X492 1 M2_M1_CDNS_765158229098 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X493 1 M2_M1_CDNS_765158229098 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X494 1 M2_M1_CDNS_765158229098 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X495 1 M2_M1_CDNS_765158229098 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X496 1 M2_M1_CDNS_765158229098 $T=30630 7680 0 0 $X=30270 $Y=7550
X497 1 M2_M1_CDNS_765158229098 $T=30630 13130 0 0 $X=30270 $Y=13000
X498 1 M9_M8_CDNS_765158229099 $T=-58270 -16370 0 0 $X=-58630 $Y=-16500
X499 1 M9_M8_CDNS_765158229099 $T=-58270 -7010 0 0 $X=-58630 $Y=-7140
X500 1 M9_M8_CDNS_765158229099 $T=-58270 4550 0 0 $X=-58630 $Y=4420
X501 1 M9_M8_CDNS_765158229099 $T=-58270 14410 0 0 $X=-58630 $Y=14280
X502 2 M9_M8_CDNS_765158229099 $T=-56610 -11840 0 0 $X=-56970 $Y=-11970
X503 2 M9_M8_CDNS_765158229099 $T=-56610 -5390 0 0 $X=-56970 $Y=-5520
X504 2 M9_M8_CDNS_765158229099 $T=-56610 9310 0 0 $X=-56970 $Y=9180
X505 2 M9_M8_CDNS_765158229099 $T=-56100 19570 0 0 $X=-56460 $Y=19440
X506 1 M9_M8_CDNS_765158229099 $T=-50900 -22240 0 0 $X=-51260 $Y=-22370
X507 1 M9_M8_CDNS_765158229099 $T=-50900 -11900 0 0 $X=-51260 $Y=-12030
X508 1 M9_M8_CDNS_765158229099 $T=-49890 -2060 0 0 $X=-50250 $Y=-2190
X509 1 M9_M8_CDNS_765158229099 $T=-49890 7690 0 0 $X=-50250 $Y=7560
X510 2 M9_M8_CDNS_765158229099 $T=-46220 -15100 0 0 $X=-46580 $Y=-15230
X511 2 M9_M8_CDNS_765158229099 $T=-46220 -6560 0 0 $X=-46580 $Y=-6690
X512 2 M9_M8_CDNS_765158229099 $T=-46220 1650 0 0 $X=-46580 $Y=1520
X513 2 M9_M8_CDNS_765158229099 $T=-46220 11880 0 0 $X=-46580 $Y=11750
X514 1 M9_M8_CDNS_765158229099 $T=-44430 -20980 0 0 $X=-44790 $Y=-21110
X515 1 M9_M8_CDNS_765158229099 $T=-44430 -12140 0 0 $X=-44790 $Y=-12270
X516 1 M9_M8_CDNS_765158229099 $T=-44430 -4800 0 0 $X=-44790 $Y=-4930
X517 1 M9_M8_CDNS_765158229099 $T=-44430 3730 0 0 $X=-44790 $Y=3600
X518 1 M9_M8_CDNS_765158229099 $T=-28700 -21260 0 0 $X=-29060 $Y=-21390
X519 1 M9_M8_CDNS_765158229099 $T=-28700 -13910 0 0 $X=-29060 $Y=-14040
X520 1 M9_M8_CDNS_765158229099 $T=-27880 -29130 0 0 $X=-28240 $Y=-29260
X521 1 M9_M8_CDNS_765158229099 $T=-25440 -5210 0 0 $X=-25800 $Y=-5340
X522 2 M9_M8_CDNS_765158229099 $T=-24070 -23850 0 0 $X=-24430 $Y=-23980
X523 2 M9_M8_CDNS_765158229099 $T=-24070 -15330 0 0 $X=-24430 $Y=-15460
X524 2 M9_M8_CDNS_765158229099 $T=-24070 -6560 0 0 $X=-24430 $Y=-6690
X525 2 M9_M8_CDNS_765158229099 $T=-24070 2480 0 0 $X=-24430 $Y=2350
X526 2 M9_M8_CDNS_765158229099 $T=-24070 21730 0 0 $X=-24430 $Y=21600
X527 1 M9_M8_CDNS_765158229099 $T=-21770 -12140 0 0 $X=-22130 $Y=-12270
X528 1 M9_M8_CDNS_765158229099 $T=-18480 -29300 0 0 $X=-18840 $Y=-29430
X529 1 M9_M8_CDNS_765158229099 $T=-18480 -21090 0 0 $X=-18840 $Y=-21220
X530 1 M9_M8_CDNS_765158229099 $T=-17260 -4900 0 0 $X=-17620 $Y=-5030
X531 1 M9_M8_CDNS_765158229099 $T=-1360 -29920 0 0 $X=-1720 $Y=-30050
X532 1 M9_M8_CDNS_765158229099 $T=-1360 -21990 0 0 $X=-1720 $Y=-22120
X533 1 M9_M8_CDNS_765158229099 $T=-1360 -14120 0 0 $X=-1720 $Y=-14250
X534 1 M9_M8_CDNS_765158229099 $T=-1190 -38350 0 0 $X=-1550 $Y=-38480
X535 2 M9_M8_CDNS_765158229099 $T=1060 -31550 0 0 $X=700 $Y=-31680
X536 2 M9_M8_CDNS_765158229099 $T=1060 -24120 0 0 $X=700 $Y=-24250
X537 2 M9_M8_CDNS_765158229099 $T=1060 -14890 0 0 $X=700 $Y=-15020
X538 2 M9_M8_CDNS_765158229099 $T=2890 -7750 0 0 $X=2530 $Y=-7880
X539 1 M9_M8_CDNS_765158229099 $T=7430 -37100 0 0 $X=7070 $Y=-37230
X540 1 M9_M8_CDNS_765158229099 $T=9050 -29250 0 0 $X=8690 $Y=-29380
X541 1 M9_M8_CDNS_765158229099 $T=9050 -19900 0 0 $X=8690 $Y=-20030
X542 1 M9_M8_CDNS_765158229099 $T=9050 -13120 0 0 $X=8690 $Y=-13250
X543 2 M9_M8_CDNS_765158229099 $T=23880 13850 0 0 $X=23520 $Y=13720
X544 2 M9_M8_CDNS_765158229099 $T=24550 3710 0 0 $X=24190 $Y=3580
X545 2 M9_M8_CDNS_765158229099 $T=26060 -34250 0 0 $X=25700 $Y=-34380
X546 2 M9_M8_CDNS_765158229099 $T=26060 -26210 0 0 $X=25700 $Y=-26340
X547 2 M9_M8_CDNS_765158229099 $T=26060 -19020 0 0 $X=25700 $Y=-19150
X548 2 M9_M8_CDNS_765158229099 $T=26060 -9950 0 0 $X=25700 $Y=-10080
X549 2 M9_M8_CDNS_765158229099 $T=29710 19070 0 0 $X=29350 $Y=18940
X550 1 M9_M8_CDNS_765158229099 $T=30630 -38350 0 0 $X=30270 $Y=-38480
X551 1 M9_M8_CDNS_765158229099 $T=30630 -29960 0 0 $X=30270 $Y=-30090
X552 1 M9_M8_CDNS_765158229099 $T=30630 -21570 0 0 $X=30270 $Y=-21700
X553 1 M9_M8_CDNS_765158229099 $T=30630 -13180 0 0 $X=30270 $Y=-13310
X554 1 M9_M8_CDNS_765158229099 $T=30630 -2200 0 0 $X=30270 $Y=-2330
X555 1 M9_M8_CDNS_765158229099 $T=30630 7680 0 0 $X=30270 $Y=7550
X556 1 M9_M8_CDNS_765158229099 $T=30630 13130 0 0 $X=30270 $Y=13000
X557 3 M5_M4_CDNS_7651582290910 $T=-32480 -13040 0 0 $X=-32560 $Y=-13170
X558 4 M5_M4_CDNS_7651582290910 $T=-31620 -4240 0 0 $X=-31700 $Y=-4370
X559 3 M5_M4_CDNS_7651582290910 $T=-31100 -13040 0 0 $X=-31180 $Y=-13170
X560 5 M5_M4_CDNS_7651582290910 $T=-30250 8200 0 0 $X=-30330 $Y=8070
X561 4 M5_M4_CDNS_7651582290910 $T=-29690 -4240 0 0 $X=-29770 $Y=-4370
X562 5 M5_M4_CDNS_7651582290910 $T=-27060 8200 0 0 $X=-27140 $Y=8070
X563 6 M5_M4_CDNS_7651582290910 $T=-6460 5940 0 0 $X=-6540 $Y=5810
X564 6 M5_M4_CDNS_7651582290910 $T=-1780 5950 0 0 $X=-1860 $Y=5820
X565 5 M2_M1_CDNS_7651582290911 $T=-62770 7460 0 0 $X=-62850 $Y=7050
X566 7 M2_M1_CDNS_7651582290911 $T=-62770 17260 0 0 $X=-62850 $Y=16850
X567 3 M2_M1_CDNS_7651582290911 $T=-62470 -13270 0 0 $X=-62550 $Y=-13680
X568 4 M2_M1_CDNS_7651582290911 $T=-62470 -3810 0 0 $X=-62550 $Y=-4220
X569 8 M2_M1_CDNS_7651582290911 $T=-61470 7170 0 0 $X=-61550 $Y=6760
X570 8 M2_M1_CDNS_7651582290911 $T=-61470 16960 0 0 $X=-61550 $Y=16550
X571 8 M2_M1_CDNS_7651582290911 $T=-61170 -13570 0 0 $X=-61250 $Y=-13980
X572 8 M2_M1_CDNS_7651582290911 $T=-61170 -4100 0 0 $X=-61250 $Y=-4510
X573 3 M2_M1_CDNS_7651582290911 $T=-54250 -18890 0 0 $X=-54330 $Y=-19300
X574 4 M2_M1_CDNS_7651582290911 $T=-54150 -8650 0 0 $X=-54230 $Y=-9060
X575 5 M2_M1_CDNS_7651582290911 $T=-54150 600 0 0 $X=-54230 $Y=190
X576 7 M2_M1_CDNS_7651582290911 $T=-54150 10410 0 0 $X=-54230 $Y=10000
X577 9 M2_M1_CDNS_7651582290911 $T=-52950 -19200 0 0 $X=-53030 $Y=-19610
X578 9 M2_M1_CDNS_7651582290911 $T=-52850 -8950 0 0 $X=-52930 $Y=-9360
X579 9 M2_M1_CDNS_7651582290911 $T=-52850 300 0 0 $X=-52930 $Y=-110
X580 9 M2_M1_CDNS_7651582290911 $T=-52850 10130 0 0 $X=-52930 $Y=9720
X581 3 M2_M1_CDNS_7651582290911 $T=-32630 -26510 0 0 $X=-32710 $Y=-26920
X582 4 M2_M1_CDNS_7651582290911 $T=-31780 -17870 0 0 $X=-31860 $Y=-18280
X583 10 M2_M1_CDNS_7651582290911 $T=-31330 -26810 0 0 $X=-31410 $Y=-27220
X584 5 M2_M1_CDNS_7651582290911 $T=-30580 -9750 0 0 $X=-30660 $Y=-10160
X585 10 M2_M1_CDNS_7651582290911 $T=-30480 -18170 0 0 $X=-30560 $Y=-18580
X586 10 M2_M1_CDNS_7651582290911 $T=-29280 -10050 0 0 $X=-29360 $Y=-10460
X587 7 M2_M1_CDNS_7651582290911 $T=-28690 -1560 0 0 $X=-28770 $Y=-1970
X588 10 M2_M1_CDNS_7651582290911 $T=-27390 -1860 0 0 $X=-27470 $Y=-2270
X589 3 M2_M1_CDNS_7651582290911 $T=-6190 -36090 0 0 $X=-6270 $Y=-36500
X590 4 M2_M1_CDNS_7651582290911 $T=-5950 -26840 0 0 $X=-6030 $Y=-27250
X591 5 M2_M1_CDNS_7651582290911 $T=-5400 -18740 0 0 $X=-5480 $Y=-19150
X592 11 M2_M1_CDNS_7651582290911 $T=-4890 -36400 0 0 $X=-4970 $Y=-36810
X593 11 M2_M1_CDNS_7651582290911 $T=-4650 -27140 0 0 $X=-4730 $Y=-27550
X594 11 M2_M1_CDNS_7651582290911 $T=-4100 -19040 0 0 $X=-4180 $Y=-19450
X595 7 M2_M1_CDNS_7651582290911 $T=-3970 -10680 0 0 $X=-4050 $Y=-11090
X596 11 M2_M1_CDNS_7651582290911 $T=-2670 -10980 0 0 $X=-2750 $Y=-11390
X597 5 M3_M2_CDNS_7651582290912 $T=-62770 7460 0 0 $X=-62850 $Y=7050
X598 7 M3_M2_CDNS_7651582290912 $T=-62770 17260 0 0 $X=-62850 $Y=16850
X599 3 M3_M2_CDNS_7651582290912 $T=-62470 -13270 0 0 $X=-62550 $Y=-13680
X600 4 M3_M2_CDNS_7651582290912 $T=-62470 -3810 0 0 $X=-62550 $Y=-4220
X601 8 M3_M2_CDNS_7651582290912 $T=-61470 7170 0 0 $X=-61550 $Y=6760
X602 8 M3_M2_CDNS_7651582290912 $T=-61470 16960 0 0 $X=-61550 $Y=16550
X603 8 M3_M2_CDNS_7651582290912 $T=-61170 -13570 0 0 $X=-61250 $Y=-13980
X604 8 M3_M2_CDNS_7651582290912 $T=-61170 -4100 0 0 $X=-61250 $Y=-4510
X605 3 M3_M2_CDNS_7651582290912 $T=-54250 -18890 0 0 $X=-54330 $Y=-19300
X606 4 M3_M2_CDNS_7651582290912 $T=-54150 -8650 0 0 $X=-54230 $Y=-9060
X607 5 M3_M2_CDNS_7651582290912 $T=-54150 600 0 0 $X=-54230 $Y=190
X608 7 M3_M2_CDNS_7651582290912 $T=-54150 10410 0 0 $X=-54230 $Y=10000
X609 9 M3_M2_CDNS_7651582290912 $T=-52950 -19200 0 0 $X=-53030 $Y=-19610
X610 9 M3_M2_CDNS_7651582290912 $T=-52850 -8950 0 0 $X=-52930 $Y=-9360
X611 9 M3_M2_CDNS_7651582290912 $T=-52850 300 0 0 $X=-52930 $Y=-110
X612 9 M3_M2_CDNS_7651582290912 $T=-52850 10130 0 0 $X=-52930 $Y=9720
X613 3 M3_M2_CDNS_7651582290912 $T=-32630 -26510 0 0 $X=-32710 $Y=-26920
X614 4 M3_M2_CDNS_7651582290912 $T=-31780 -17870 0 0 $X=-31860 $Y=-18280
X615 10 M3_M2_CDNS_7651582290912 $T=-31330 -26810 0 0 $X=-31410 $Y=-27220
X616 5 M3_M2_CDNS_7651582290912 $T=-30580 -9750 0 0 $X=-30660 $Y=-10160
X617 10 M3_M2_CDNS_7651582290912 $T=-30480 -18170 0 0 $X=-30560 $Y=-18580
X618 10 M3_M2_CDNS_7651582290912 $T=-29280 -10050 0 0 $X=-29360 $Y=-10460
X619 7 M3_M2_CDNS_7651582290912 $T=-28690 -1560 0 0 $X=-28770 $Y=-1970
X620 10 M3_M2_CDNS_7651582290912 $T=-27390 -1860 0 0 $X=-27470 $Y=-2270
X621 3 M3_M2_CDNS_7651582290912 $T=-6190 -36090 0 0 $X=-6270 $Y=-36500
X622 4 M3_M2_CDNS_7651582290912 $T=-5950 -26840 0 0 $X=-6030 $Y=-27250
X623 5 M3_M2_CDNS_7651582290912 $T=-5400 -18740 0 0 $X=-5480 $Y=-19150
X624 11 M3_M2_CDNS_7651582290912 $T=-4890 -36400 0 0 $X=-4970 $Y=-36810
X625 11 M3_M2_CDNS_7651582290912 $T=-4650 -27140 0 0 $X=-4730 $Y=-27550
X626 11 M3_M2_CDNS_7651582290912 $T=-4100 -19040 0 0 $X=-4180 $Y=-19450
X627 7 M3_M2_CDNS_7651582290912 $T=-3970 -10680 0 0 $X=-4050 $Y=-11090
X628 11 M3_M2_CDNS_7651582290912 $T=-2670 -10980 0 0 $X=-2750 $Y=-11390
X629 5 M4_M3_CDNS_7651582290913 $T=-62770 7460 0 0 $X=-62850 $Y=7050
X630 7 M4_M3_CDNS_7651582290913 $T=-62770 17260 0 0 $X=-62850 $Y=16850
X631 3 M4_M3_CDNS_7651582290913 $T=-62470 -13270 0 0 $X=-62550 $Y=-13680
X632 4 M4_M3_CDNS_7651582290913 $T=-62470 -3810 0 0 $X=-62550 $Y=-4220
X633 3 M4_M3_CDNS_7651582290913 $T=-54250 -18890 0 0 $X=-54330 $Y=-19300
X634 7 M4_M3_CDNS_7651582290913 $T=-54160 10400 0 0 $X=-54240 $Y=9990
X635 4 M4_M3_CDNS_7651582290913 $T=-54150 -8650 0 0 $X=-54230 $Y=-9060
X636 5 M4_M3_CDNS_7651582290913 $T=-54150 600 0 0 $X=-54230 $Y=190
X637 3 M4_M3_CDNS_7651582290913 $T=-32630 -26510 0 0 $X=-32710 $Y=-26920
X638 4 M4_M3_CDNS_7651582290913 $T=-31780 -17870 0 0 $X=-31860 $Y=-18280
X639 5 M4_M3_CDNS_7651582290913 $T=-30580 -9750 0 0 $X=-30660 $Y=-10160
X640 7 M4_M3_CDNS_7651582290913 $T=-28690 -1560 0 0 $X=-28770 $Y=-1970
X641 3 M4_M3_CDNS_7651582290913 $T=-6190 -36090 0 0 $X=-6270 $Y=-36500
X642 4 M4_M3_CDNS_7651582290913 $T=-5950 -26840 0 0 $X=-6030 $Y=-27250
X643 5 M4_M3_CDNS_7651582290913 $T=-5400 -18740 0 0 $X=-5480 $Y=-19150
X644 7 M4_M3_CDNS_7651582290913 $T=-3970 -10680 0 0 $X=-4050 $Y=-11090
X645 12 M2_M1_CDNS_7651582290914 $T=-59460 7520 0 0 $X=-59540 $Y=7390
X646 13 M2_M1_CDNS_7651582290914 $T=-59450 17310 0 0 $X=-59530 $Y=17180
X647 14 M2_M1_CDNS_7651582290914 $T=-59160 -13210 0 0 $X=-59240 $Y=-13340
X648 15 M2_M1_CDNS_7651582290914 $T=-59160 -3740 0 0 $X=-59240 $Y=-3870
X649 16 M2_M1_CDNS_7651582290914 $T=-50940 -18840 0 0 $X=-51020 $Y=-18970
X650 17 M2_M1_CDNS_7651582290914 $T=-50840 650 0 0 $X=-50920 $Y=520
X651 18 M2_M1_CDNS_7651582290914 $T=-50840 10480 0 0 $X=-50920 $Y=10350
X652 19 M2_M1_CDNS_7651582290914 $T=-50830 -8590 0 0 $X=-50910 $Y=-8720
X653 20 M2_M1_CDNS_7651582290914 $T=-29320 -26450 0 0 $X=-29400 $Y=-26580
X654 21 M2_M1_CDNS_7651582290914 $T=-28460 -17820 0 0 $X=-28540 $Y=-17950
X655 22 M2_M1_CDNS_7651582290914 $T=-27220 -9690 0 0 $X=-27300 $Y=-9820
X656 23 M2_M1_CDNS_7651582290914 $T=-25370 -1500 0 0 $X=-25450 $Y=-1630
X657 24 M2_M1_CDNS_7651582290914 $T=-2890 -36050 0 0 $X=-2970 $Y=-36180
X658 25 M2_M1_CDNS_7651582290914 $T=-2630 -26770 0 0 $X=-2710 $Y=-26900
X659 26 M2_M1_CDNS_7651582290914 $T=-2090 -18700 0 0 $X=-2170 $Y=-18830
X660 27 M2_M1_CDNS_7651582290914 $T=-660 -10620 0 0 $X=-740 $Y=-10750
X661 24 M2_M1_CDNS_7651582290914 $T=8560 -32030 0 0 $X=8480 $Y=-32160
X662 25 M2_M1_CDNS_7651582290914 $T=8560 -24560 0 0 $X=8480 $Y=-24690
X663 26 M2_M1_CDNS_7651582290914 $T=8560 -15380 0 0 $X=8480 $Y=-15510
X664 27 M2_M1_CDNS_7651582290914 $T=8560 -8150 0 0 $X=8480 $Y=-8280
X665 28 M2_M1_CDNS_7651582290914 $T=18160 -35920 0 0 $X=18080 $Y=-36050
X666 29 M2_M1_CDNS_7651582290914 $T=18160 -28450 0 0 $X=18080 $Y=-28580
X667 30 M2_M1_CDNS_7651582290914 $T=18160 -19270 0 0 $X=18080 $Y=-19400
X668 31 M2_M1_CDNS_7651582290914 $T=18160 -12040 0 0 $X=18080 $Y=-12170
X669 32 M2_M1_CDNS_7651582290914 $T=24420 1860 0 0 $X=24340 $Y=1730
X670 6 M2_M1_CDNS_7651582290914 $T=24420 11860 0 0 $X=24340 $Y=11730
X671 13 M2_M1_CDNS_7651582290914 $T=29830 17270 0 0 $X=29750 $Y=17140
X672 16 M3_M2_CDNS_7651582290915 $T=-50940 -18840 0 0 $X=-51020 $Y=-18970
X673 33 M3_M2_CDNS_7651582290915 $T=-47750 -8680 0 0 $X=-47830 $Y=-8810
X674 34 M3_M2_CDNS_7651582290915 $T=-47550 -600 0 0 $X=-47630 $Y=-730
X675 19 M3_M2_CDNS_7651582290915 $T=-47140 -9690 0 0 $X=-47220 $Y=-9820
X676 14 M3_M2_CDNS_7651582290915 $T=-47100 -10630 0 0 $X=-47180 $Y=-10760
X677 15 M3_M2_CDNS_7651582290915 $T=-46210 -2290 0 0 $X=-46290 $Y=-2420
X678 17 M3_M2_CDNS_7651582290915 $T=-46200 -1350 0 0 $X=-46280 $Y=-1480
X679 35 M3_M2_CDNS_7651582290915 $T=-45000 -17050 0 0 $X=-45080 $Y=-17180
X680 18 M3_M2_CDNS_7651582290915 $T=-43770 6810 0 0 $X=-43850 $Y=6680
X681 12 M3_M2_CDNS_7651582290915 $T=-43760 6340 0 0 $X=-43840 $Y=6210
X682 21 M3_M2_CDNS_7651582290915 $T=-26920 -17820 0 0 $X=-27000 $Y=-17950
X683 20 M3_M2_CDNS_7651582290915 $T=-26910 -26460 0 0 $X=-26990 $Y=-26590
X684 36 M3_M2_CDNS_7651582290915 $T=-25730 -27040 0 0 $X=-25810 $Y=-27170
X685 22 M3_M2_CDNS_7651582290915 $T=-25010 -9690 0 0 $X=-25090 $Y=-9820
X686 23 M3_M2_CDNS_7651582290915 $T=-23170 -1500 0 0 $X=-23250 $Y=-1630
X687 37 M3_M2_CDNS_7651582290915 $T=-22130 -18280 0 0 $X=-22210 $Y=-18410
X688 38 M3_M2_CDNS_7651582290915 $T=-22050 -10130 0 0 $X=-22130 $Y=-10260
X689 39 M3_M2_CDNS_7651582290915 $T=-22000 -26530 0 0 $X=-22080 $Y=-26660
X690 25 M3_M2_CDNS_7651582290915 $T=-140 -26730 0 0 $X=-220 $Y=-26860
X691 24 M3_M2_CDNS_7651582290915 $T=50 -35270 0 0 $X=-30 $Y=-35400
X692 26 M3_M2_CDNS_7651582290915 $T=200 -18330 0 0 $X=120 $Y=-18460
X693 24 M3_M2_CDNS_7651582290915 $T=7210 -32030 0 0 $X=7130 $Y=-32160
X694 25 M3_M2_CDNS_7651582290915 $T=7210 -24560 0 0 $X=7130 $Y=-24690
X695 26 M3_M2_CDNS_7651582290915 $T=7210 -15380 0 0 $X=7130 $Y=-15510
X696 29 M3_M2_CDNS_7651582290915 $T=16810 -28450 0 0 $X=16730 $Y=-28580
X697 30 M3_M2_CDNS_7651582290915 $T=16810 -19270 0 0 $X=16730 $Y=-19400
X698 31 M3_M2_CDNS_7651582290915 $T=16810 -12040 0 0 $X=16730 $Y=-12170
X699 32 M3_M2_CDNS_7651582290915 $T=23070 1860 0 0 $X=22990 $Y=1730
X700 6 M3_M2_CDNS_7651582290915 $T=23070 11860 0 0 $X=22990 $Y=11730
X701 40 M3_M2_CDNS_7651582290915 $T=28730 -18680 0 0 $X=28650 $Y=-18810
X702 41 M3_M2_CDNS_7651582290915 $T=28820 -35530 0 0 $X=28740 $Y=-35660
X703 42 M3_M2_CDNS_7651582290915 $T=29100 -27090 0 0 $X=29020 $Y=-27220
X704 43 M2_M1_CDNS_7651582290916 $T=15160 -33790 0 0 $X=14940 $Y=-33920
X705 43 M2_M1_CDNS_7651582290916 $T=15160 -26320 0 0 $X=14940 $Y=-26450
X706 43 M2_M1_CDNS_7651582290916 $T=15160 -17140 0 0 $X=14940 $Y=-17270
X707 43 M2_M1_CDNS_7651582290916 $T=15160 -9950 0 0 $X=14940 $Y=-10080
X708 44 M2_M1_CDNS_7651582290916 $T=16040 -32690 0 0 $X=15820 $Y=-32820
X709 45 M2_M1_CDNS_7651582290916 $T=16040 -25220 0 0 $X=15820 $Y=-25350
X710 46 M2_M1_CDNS_7651582290916 $T=16040 -16040 0 0 $X=15820 $Y=-16170
X711 47 M2_M1_CDNS_7651582290916 $T=16040 -8810 0 0 $X=15820 $Y=-8940
X712 43 M2_M1_CDNS_7651582290916 $T=24760 -37680 0 0 $X=24540 $Y=-37810
X713 43 M2_M1_CDNS_7651582290916 $T=24760 -30210 0 0 $X=24540 $Y=-30340
X714 43 M2_M1_CDNS_7651582290916 $T=24760 -21030 0 0 $X=24540 $Y=-21160
X715 43 M2_M1_CDNS_7651582290916 $T=24760 -13800 0 0 $X=24540 $Y=-13930
X716 48 M2_M1_CDNS_7651582290916 $T=25640 -36580 0 0 $X=25420 $Y=-36710
X717 49 M2_M1_CDNS_7651582290916 $T=25640 -29110 0 0 $X=25420 $Y=-29240
X718 50 M2_M1_CDNS_7651582290916 $T=25640 -19930 0 0 $X=25420 $Y=-20060
X719 51 M2_M1_CDNS_7651582290916 $T=25640 -12700 0 0 $X=25420 $Y=-12830
X720 43 M2_M1_CDNS_7651582290916 $T=30980 10090 0 0 $X=30760 $Y=9960
X721 43 M2_M1_CDNS_7651582290916 $T=31010 50 0 0 $X=30790 $Y=-80
X722 52 M2_M1_CDNS_7651582290916 $T=31900 1200 0 0 $X=31680 $Y=1070
X723 53 M2_M1_CDNS_7651582290916 $T=31900 11200 0 0 $X=31680 $Y=11070
X724 43 M2_M1_CDNS_7651582290916 $T=36420 15480 0 0 $X=36200 $Y=15350
X725 54 M2_M1_CDNS_7651582290916 $T=37310 16610 0 0 $X=37090 $Y=16480
X726 55 M4_M3_CDNS_7651582290917 $T=7590 -25970 0 0 $X=7370 $Y=-26100
X727 55 M4_M3_CDNS_7651582290917 $T=7590 -16790 0 0 $X=7370 $Y=-16920
X728 55 M4_M3_CDNS_7651582290917 $T=7590 -9560 0 0 $X=7370 $Y=-9690
X729 55 M4_M3_CDNS_7651582290917 $T=7600 -33440 0 0 $X=7380 $Y=-33570
X730 43 M4_M3_CDNS_7651582290917 $T=15160 -33790 0 0 $X=14940 $Y=-33920
X731 43 M4_M3_CDNS_7651582290917 $T=15160 -26320 0 0 $X=14940 $Y=-26450
X732 43 M4_M3_CDNS_7651582290917 $T=15160 -17140 0 0 $X=14940 $Y=-17270
X733 43 M4_M3_CDNS_7651582290917 $T=15160 -9950 0 0 $X=14940 $Y=-10080
X734 55 M4_M3_CDNS_7651582290917 $T=17180 -5650 0 0 $X=16960 $Y=-5780
X735 55 M4_M3_CDNS_7651582290917 $T=17180 -3660 0 0 $X=16960 $Y=-3790
X736 55 M4_M3_CDNS_7651582290917 $T=17190 -37330 0 0 $X=16970 $Y=-37460
X737 55 M4_M3_CDNS_7651582290917 $T=17190 -29860 0 0 $X=16970 $Y=-29990
X738 55 M4_M3_CDNS_7651582290917 $T=17190 -20680 0 0 $X=16970 $Y=-20810
X739 55 M4_M3_CDNS_7651582290917 $T=17190 -13450 0 0 $X=16970 $Y=-13580
X740 55 M4_M3_CDNS_7651582290917 $T=23440 10450 0 0 $X=23220 $Y=10320
X741 55 M4_M3_CDNS_7651582290917 $T=23450 450 0 0 $X=23230 $Y=320
X742 43 M4_M3_CDNS_7651582290917 $T=24760 -37680 0 180 $X=24540 $Y=-37810
X743 43 M4_M3_CDNS_7651582290917 $T=24760 -30210 0 180 $X=24540 $Y=-30340
X744 43 M4_M3_CDNS_7651582290917 $T=24760 -21030 0 180 $X=24540 $Y=-21160
X745 43 M4_M3_CDNS_7651582290917 $T=24760 -13800 0 0 $X=24540 $Y=-13930
X746 55 M4_M3_CDNS_7651582290917 $T=25000 20350 0 0 $X=24780 $Y=20220
X747 55 M4_M3_CDNS_7651582290917 $T=28860 15860 0 0 $X=28640 $Y=15730
X748 43 M4_M3_CDNS_7651582290917 $T=30980 10090 0 0 $X=30760 $Y=9960
X749 43 M4_M3_CDNS_7651582290917 $T=31010 50 0 0 $X=30790 $Y=-80
X750 43 M4_M3_CDNS_7651582290917 $T=36420 15480 0 0 $X=36200 $Y=15350
X751 43 M4_M3_CDNS_7651582290917 $T=36420 20180 0 0 $X=36200 $Y=20050
X752 55 M3_M2_CDNS_7651582290918 $T=7590 -33440 0 0 $X=7370 $Y=-33570
X753 55 M3_M2_CDNS_7651582290918 $T=7590 -25970 0 0 $X=7370 $Y=-26100
X754 55 M3_M2_CDNS_7651582290918 $T=7590 -16790 0 0 $X=7370 $Y=-16920
X755 55 M3_M2_CDNS_7651582290918 $T=7590 -9560 0 0 $X=7370 $Y=-9690
X756 43 M3_M2_CDNS_7651582290918 $T=15160 -33790 0 0 $X=14940 $Y=-33920
X757 43 M3_M2_CDNS_7651582290918 $T=15160 -26320 0 0 $X=14940 $Y=-26450
X758 43 M3_M2_CDNS_7651582290918 $T=15160 -17140 0 0 $X=14940 $Y=-17270
X759 43 M3_M2_CDNS_7651582290918 $T=15160 -9950 0 0 $X=14940 $Y=-10080
X760 44 M3_M2_CDNS_7651582290918 $T=16040 -32690 0 0 $X=15820 $Y=-32820
X761 45 M3_M2_CDNS_7651582290918 $T=16040 -25220 0 0 $X=15820 $Y=-25350
X762 46 M3_M2_CDNS_7651582290918 $T=16040 -16040 0 0 $X=15820 $Y=-16170
X763 47 M3_M2_CDNS_7651582290918 $T=16040 -8810 0 0 $X=15820 $Y=-8940
X764 55 M3_M2_CDNS_7651582290918 $T=17190 -37330 0 0 $X=16970 $Y=-37460
X765 55 M3_M2_CDNS_7651582290918 $T=17190 -29860 0 0 $X=16970 $Y=-29990
X766 55 M3_M2_CDNS_7651582290918 $T=17190 -20680 0 0 $X=16970 $Y=-20810
X767 55 M3_M2_CDNS_7651582290918 $T=17190 -13450 0 0 $X=16970 $Y=-13580
X768 55 M3_M2_CDNS_7651582290918 $T=23450 450 0 0 $X=23230 $Y=320
X769 55 M3_M2_CDNS_7651582290918 $T=23450 10450 0 0 $X=23230 $Y=10320
X770 43 M3_M2_CDNS_7651582290918 $T=24760 -37680 0 0 $X=24540 $Y=-37810
X771 43 M3_M2_CDNS_7651582290918 $T=24760 -30210 0 0 $X=24540 $Y=-30340
X772 43 M3_M2_CDNS_7651582290918 $T=24760 -21030 0 0 $X=24540 $Y=-21160
X773 43 M3_M2_CDNS_7651582290918 $T=24760 -13800 0 0 $X=24540 $Y=-13930
X774 48 M3_M2_CDNS_7651582290918 $T=25640 -36580 0 0 $X=25420 $Y=-36710
X775 49 M3_M2_CDNS_7651582290918 $T=25640 -29110 0 0 $X=25420 $Y=-29240
X776 50 M3_M2_CDNS_7651582290918 $T=25640 -19930 0 0 $X=25420 $Y=-20060
X777 51 M3_M2_CDNS_7651582290918 $T=25640 -12700 0 0 $X=25420 $Y=-12830
X778 55 M3_M2_CDNS_7651582290918 $T=28860 15860 0 0 $X=28640 $Y=15730
X779 43 M3_M2_CDNS_7651582290918 $T=30980 10090 0 0 $X=30760 $Y=9960
X780 43 M3_M2_CDNS_7651582290918 $T=31010 50 0 0 $X=30790 $Y=-80
X781 52 M3_M2_CDNS_7651582290918 $T=31900 1200 0 0 $X=31680 $Y=1070
X782 53 M3_M2_CDNS_7651582290918 $T=31900 11200 0 0 $X=31680 $Y=11070
X783 43 M3_M2_CDNS_7651582290918 $T=36420 15480 0 0 $X=36200 $Y=15350
X784 54 M3_M2_CDNS_7651582290918 $T=37310 16610 0 0 $X=37090 $Y=16480
X785 56 M4_M3_CDNS_7651582290919 $T=-31890 -19910 0 0 $X=-31970 $Y=-20040
X786 57 M4_M3_CDNS_7651582290919 $T=-31130 -10620 0 0 $X=-31210 $Y=-10750
X787 58 M4_M3_CDNS_7651582290919 $T=-29610 -3090 0 0 $X=-29690 $Y=-3220
X788 6 M4_M3_CDNS_7651582290919 $T=-28160 5940 0 0 $X=-28240 $Y=5810
X789 56 M4_M3_CDNS_7651582290919 $T=-27090 -19910 0 0 $X=-27170 $Y=-20040
X790 57 M4_M3_CDNS_7651582290919 $T=-26310 -10630 0 0 $X=-26390 $Y=-10760
X791 58 M4_M3_CDNS_7651582290919 $T=-23220 -3090 0 0 $X=-23300 $Y=-3220
X792 29 M4_M3_CDNS_7651582290919 $T=-5630 -29010 0 0 $X=-5710 $Y=-29140
X793 30 M4_M3_CDNS_7651582290919 $T=-5420 -20630 0 0 $X=-5500 $Y=-20760
X794 31 M4_M3_CDNS_7651582290919 $T=-4530 -12400 0 0 $X=-4610 $Y=-12530
X795 32 M4_M3_CDNS_7651582290919 $T=-3390 -2610 0 0 $X=-3470 $Y=-2740
X796 29 M4_M3_CDNS_7651582290919 $T=-1190 -29010 0 0 $X=-1270 $Y=-29140
X797 30 M4_M3_CDNS_7651582290919 $T=-50 -20630 0 0 $X=-130 $Y=-20760
X798 31 M4_M3_CDNS_7651582290919 $T=890 -12410 0 0 $X=810 $Y=-12540
X799 32 M4_M3_CDNS_7651582290919 $T=20010 1820 0 0 $X=19930 $Y=1690
X800 6 M4_M3_CDNS_7651582290919 $T=20870 11820 0 0 $X=20790 $Y=11690
X801 3 M4_M3_CDNS_7651582290920 $T=-65780 -13030 0 0 $X=-66140 $Y=-13520
X802 4 M4_M3_CDNS_7651582290920 $T=-65680 -4250 0 0 $X=-66040 $Y=-4740
X803 5 M4_M3_CDNS_7651582290921 $T=-65760 8200 0 0 $X=-66200 $Y=7790
X804 7 M4_M3_CDNS_7651582290921 $T=-65570 17450 0 0 $X=-66010 $Y=17040
X805 5 2 8 1 12 142 64 and2 $T=-60420 7100 0 0 $X=-63090 $Y=4520
X806 7 2 8 1 13 143 65 and2 $T=-60420 16900 0 0 $X=-63090 $Y=14320
X807 3 2 8 1 14 144 66 and2 $T=-60120 -13630 0 0 $X=-62790 $Y=-16210
X808 4 2 8 1 15 145 67 and2 $T=-60120 -4160 0 0 $X=-62790 $Y=-6740
X809 3 2 9 1 16 146 68 and2 $T=-51900 -19260 0 0 $X=-54570 $Y=-21840
X810 4 2 9 1 19 147 69 and2 $T=-51800 -9010 0 0 $X=-54470 $Y=-11590
X811 5 2 9 1 17 148 70 and2 $T=-51800 240 0 0 $X=-54470 $Y=-2340
X812 7 2 9 1 18 149 71 and2 $T=-51800 10060 0 0 $X=-54470 $Y=7480
X813 3 2 10 1 20 150 72 and2 $T=-30280 -26870 0 0 $X=-32950 $Y=-29450
X814 4 2 10 1 21 151 73 and2 $T=-29430 -18230 0 0 $X=-32100 $Y=-20810
X815 5 2 10 1 22 152 74 and2 $T=-28230 -10110 0 0 $X=-30900 $Y=-12690
X816 7 2 10 1 23 153 75 and2 $T=-26340 -1920 0 0 $X=-29010 $Y=-4500
X817 3 2 11 1 24 154 76 and2 $T=-3840 -36460 0 0 $X=-6510 $Y=-39040
X818 4 2 11 1 25 155 77 and2 $T=-3600 -27200 0 0 $X=-6270 $Y=-29780
X819 5 2 11 1 26 156 78 and2 $T=-3050 -19100 0 0 $X=-5720 $Y=-21680
X820 7 2 11 1 27 157 79 and2 $T=-1620 -11040 0 0 $X=-4290 $Y=-13620
X821 35 16 1 2 56 36 80 half_adder $T=-46360 -21200 0 0 $X=-44060 $Y=-20920
X822 18 12 1 2 6 34 82 half_adder $T=-46060 3240 0 0 $X=-43760 $Y=3520
X823 23 58 1 2 32 38 84 half_adder $T=-20950 -5320 0 0 $X=-18650 $Y=-5040
X824 47 51 1 2 59 40 86 half_adder $T=28740 -13320 0 0 $X=31040 $Y=-13040
X825 19 14 33 2 1 57 35 90 89 91
+ 88 full_adder $T=-47430 -13530 0 0 $X=-45650 $Y=-12280
X826 17 15 34 2 1 58 33 94 93 95
+ 92 full_adder $T=-47430 -5190 0 0 $X=-45650 $Y=-3940
X827 21 56 37 2 1 30 39 98 97 99
+ 96 full_adder $T=-22320 -21750 0 0 $X=-20540 $Y=-20500
X828 22 57 38 2 1 31 37 102 101 103
+ 100 full_adder $T=-22320 -13530 0 0 $X=-20540 $Y=-12280
X829 20 36 39 2 1 29 28 106 105 107
+ 104 full_adder $T=-21720 -29970 0 0 $X=-19940 $Y=-28720
X830 46 50 40 2 1 60 42 110 109 111
+ 108 full_adder $T=28360 -22090 0 0 $X=30140 $Y=-20840
X831 45 49 42 2 1 61 41 114 113 115
+ 112 full_adder $T=29020 -30550 0 0 $X=30800 $Y=-29300
X832 44 48 41 2 1 62 63 118 117 119
+ 116 full_adder $T=29030 -39000 0 0 $X=30810 $Y=-37750
X833 55 2 1 24 44 43 120 121 178 179 c2mos $T=7070 -35410 0 0 $X=7070 $Y=-35560
X834 55 2 1 25 45 43 122 123 180 181 c2mos $T=7070 -27940 0 0 $X=7070 $Y=-28090
X835 55 2 1 26 46 43 124 125 182 183 c2mos $T=7070 -18760 0 0 $X=7070 $Y=-18910
X836 55 2 1 27 47 43 126 127 184 185 c2mos $T=7070 -11530 0 0 $X=7070 $Y=-11680
X837 55 2 1 28 48 43 128 129 186 187 c2mos $T=16670 -39300 0 0 $X=16670 $Y=-39450
X838 55 2 1 29 49 43 130 131 188 189 c2mos $T=16670 -31830 0 0 $X=16670 $Y=-31980
X839 55 2 1 30 50 43 132 133 190 191 c2mos $T=16670 -22650 0 0 $X=16670 $Y=-22800
X840 55 2 1 31 51 43 134 135 192 193 c2mos $T=16670 -15420 0 0 $X=16670 $Y=-15570
X841 55 2 1 6 53 43 136 137 194 195 c2mos $T=22890 8490 0 0 $X=22890 $Y=8340
X842 55 2 1 32 52 43 138 139 196 197 c2mos $T=22920 -1540 0 0 $X=22920 $Y=-1690
X843 55 2 1 13 54 43 140 141 198 199 c2mos $T=28330 13890 0 0 $X=28330 $Y=13740
M0 120 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=7820 $Y=-34760 $dt=0
M1 122 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=7820 $Y=-27290 $dt=0
M2 124 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=7820 $Y=-18110 $dt=0
M3 126 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=7820 $Y=-10880 $dt=0
M4 1 43 44 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=15280 $Y=-35240 $dt=0
M5 1 43 45 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=15280 $Y=-27770 $dt=0
M6 1 43 46 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=15280 $Y=-18590 $dt=0
M7 1 43 47 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.42231 scb=0.000192056 scc=1.27713e-07 $X=15280 $Y=-11360 $dt=0
M8 128 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=17420 $Y=-38650 $dt=0
M9 130 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=17420 $Y=-31180 $dt=0
M10 132 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=17420 $Y=-22000 $dt=0
M11 134 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=17420 $Y=-14770 $dt=0
M12 136 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=23640 $Y=9140 $dt=0
M13 138 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.37831 scb=0.00150412 scc=4.69705e-06 $X=23670 $Y=-890 $dt=0
M14 1 43 48 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=24880 $Y=-39130 $dt=0
M15 1 43 49 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=24880 $Y=-31660 $dt=0
M16 1 43 50 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=24880 $Y=-22480 $dt=0
M17 1 43 51 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=24880 $Y=-15250 $dt=0
M18 140 55 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=5.48209 scb=0.00151892 scc=4.69814e-06 $X=29080 $Y=14540 $dt=0
M19 1 43 53 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=31100 $Y=8660 $dt=0
M20 1 43 52 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=31130 $Y=-1370 $dt=0
M21 1 43 54 1 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=3.26523 scb=9.5203e-05 scc=3.22105e-09 $X=36540 $Y=14060 $dt=0
M22 64 5 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-62670 $Y=8030 $dt=1
M23 65 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-62670 $Y=17830 $dt=1
M24 66 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-62370 $Y=-12700 $dt=1
M25 67 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-62370 $Y=-3230 $dt=1
M26 2 5 64 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-62260 $Y=8030 $dt=1
M27 2 7 65 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-62260 $Y=17830 $dt=1
M28 2 3 66 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-61960 $Y=-12700 $dt=1
M29 2 4 67 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-61960 $Y=-3230 $dt=1
M30 64 8 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-61370 $Y=8030 $dt=1
M31 65 8 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-61370 $Y=17830 $dt=1
M32 66 8 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-61070 $Y=-12700 $dt=1
M33 67 8 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-61070 $Y=-3230 $dt=1
M34 68 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-54150 $Y=-18330 $dt=1
M35 69 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-54050 $Y=-8080 $dt=1
M36 70 5 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-54050 $Y=1170 $dt=1
M37 71 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-54050 $Y=10990 $dt=1
M38 2 3 68 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-53740 $Y=-18330 $dt=1
M39 2 4 69 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-53640 $Y=-8080 $dt=1
M40 2 5 70 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-53640 $Y=1170 $dt=1
M41 2 7 71 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-53640 $Y=10990 $dt=1
M42 68 9 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-52850 $Y=-18330 $dt=1
M43 69 9 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-52750 $Y=-8080 $dt=1
M44 70 9 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-52750 $Y=1170 $dt=1
M45 71 9 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-52750 $Y=10990 $dt=1
M46 72 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-32530 $Y=-25940 $dt=1
M47 2 3 72 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-32120 $Y=-25940 $dt=1
M48 73 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-31680 $Y=-17300 $dt=1
M49 2 4 73 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-31270 $Y=-17300 $dt=1
M50 72 10 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-31230 $Y=-25940 $dt=1
M51 74 5 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-30480 $Y=-9180 $dt=1
M52 73 10 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-30380 $Y=-17300 $dt=1
M53 2 5 74 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-30070 $Y=-9180 $dt=1
M54 74 10 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-29180 $Y=-9180 $dt=1
M55 75 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-28590 $Y=-990 $dt=1
M56 2 7 75 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-28180 $Y=-990 $dt=1
M57 75 10 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-27290 $Y=-990 $dt=1
M58 76 3 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-6090 $Y=-35530 $dt=1
M59 77 4 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-5850 $Y=-26270 $dt=1
M60 2 3 76 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-5680 $Y=-35530 $dt=1
M61 2 4 77 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-5440 $Y=-26270 $dt=1
M62 78 5 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-5300 $Y=-18170 $dt=1
M63 2 5 78 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-4890 $Y=-18170 $dt=1
M64 76 11 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-4790 $Y=-35530 $dt=1
M65 77 11 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-4550 $Y=-26270 $dt=1
M66 78 11 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-4000 $Y=-18170 $dt=1
M67 79 7 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=-3870 $Y=-10110 $dt=1
M68 2 7 79 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=-3460 $Y=-10110 $dt=1
M69 79 11 2 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=-2570 $Y=-10110 $dt=1
.ends pipeline_mult_debug
