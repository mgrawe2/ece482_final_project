* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : xor                                          *
* Netlisted  : Sat Nov 29 12:39:47 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764441582630                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764441582630 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764441582630

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764441582631                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764441582631 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764441582631

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764441582630                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764441582630 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3034 scb=0.0125586 scc=0.000527096 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764441582630

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764441582631                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764441582631 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=39.9325 scb=0.0377946 scc=0.00385132 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764441582631

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
** N=4 EP=4 FDC=2
X0 4 2 1 nmos1v_CDNS_764441582630 $T=-50 -540 0 0 $X=-470 $Y=-740
X1 3 2 1 4 3 pmos1v_CDNS_764441582631 $T=-50 460 0 0 $X=-470 $Y=260
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764441582632                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764441582632 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=48.7608 scb=0.0470044 scc=0.00589085 $X=0 $Y=0 $dt=1
M1 3 1 2 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=56.1562 scb=0.0589139 scc=0.00666125 $X=410 $Y=0 $dt=1
.ends pmos1v_CDNS_764441582632

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764441582633                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764441582633 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=5.12155 scb=0.00103813 scc=1.48881e-06 $X=0 $Y=0 $dt=0
M1 3 1 2 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=5.12155 scb=0.00103813 scc=1.48881e-06 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764441582633

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 3 2 6 4 5
** N=6 EP=6 FDC=6
X0 1 M2_M1_CDNS_764441582630 $T=360 650 0 0 $X=280 $Y=240
X1 1 M2_M1_CDNS_764441582630 $T=1260 650 0 0 $X=1180 $Y=240
X2 2 M1_PO_CDNS_764441582631 $T=850 -1090 0 0 $X=750 $Y=-1450
X3 3 M1_PO_CDNS_764441582631 $T=850 2390 0 0 $X=750 $Y=2030
X4 1 M1_PO_CDNS_764441582631 $T=1260 650 0 0 $X=1160 $Y=290
X5 3 2 4 5 inv $T=-790 -50 0 0 $X=-1590 $Y=-1230
X6 1 6 3 5 4 pmos1v_CDNS_764441582632 $T=660 1350 0 0 $X=240 $Y=1150
X7 1 6 2 5 nmos1v_CDNS_764441582633 $T=660 -340 0 0 $X=240 $Y=-540
.ends xor
