* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : full_adder_auto                              *
* Netlisted  : Thu Dec  4 16:49:55 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888589640                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888589640 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888589640

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888589641                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888589641 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888589641

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764888589642                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764888589642 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764888589642

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888589643                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888589643 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888589643

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764888589644                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764888589644 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764888589644

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_764888589645                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_764888589645 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_764888589645

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_7648885896412                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_7648885896412 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_7648885896412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7648885896413                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7648885896413 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7648885896413

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_7648885896414                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_7648885896414 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_7648885896414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764888589640                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764888589640 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=0
.ends pmos1v_CDNS_764888589640

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764888589641                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764888589641 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 2 3 1 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 3 2 5 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
.ends nmos1v_CDNS_764888589641

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
X0 2 M1_NWELL_CDNS_7648885896412 $T=190 2570 0 0 $X=-230 $Y=2270
X1 1 M1_PO_CDNS_7648885896413 $T=-160 30 0 0 $X=-260 $Y=-330
X2 4 M1_PSUB_CDNS_7648885896414 $T=190 -2020 0 0 $X=-190 $Y=-2160
X3 2 3 1 2 4 2 pmos1v_CDNS_764888589640 $T=-60 630 0 0 $X=-480 $Y=430
X4 4 3 1 4 4 nmos1v_CDNS_764888589641 $T=-60 -1520 0 0 $X=-480 $Y=-1720
.ends inv

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764888589647                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764888589647 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764888589647

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764888589649                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764888589649 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764888589649

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xor                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xor 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=9
X0 6 M2_M1_CDNS_764888589640 $T=-30 -450 0 0 $X=-160 $Y=-580
X1 5 M2_M1_CDNS_764888589640 $T=1330 -190 0 0 $X=1200 $Y=-320
X2 6 M2_M1_CDNS_764888589641 $T=-300 -1260 0 0 $X=-430 $Y=-1390
X3 6 M2_M1_CDNS_764888589641 $T=-250 380 0 0 $X=-380 $Y=250
X4 5 M2_M1_CDNS_764888589647 $T=-660 -1560 0 0 $X=-740 $Y=-1810
X5 5 M2_M1_CDNS_764888589647 $T=-660 950 0 0 $X=-740 $Y=700
X6 5 M2_M1_CDNS_764888589647 $T=160 -1560 0 0 $X=80 $Y=-1810
X7 5 M2_M1_CDNS_764888589647 $T=160 950 0 0 $X=80 $Y=700
X8 5 M2_M1_CDNS_764888589647 $T=1050 -1560 0 0 $X=970 $Y=-1810
X9 5 M2_M1_CDNS_764888589647 $T=1050 950 0 0 $X=970 $Y=700
X10 1 M1_PO_CDNS_764888589649 $T=-450 10 0 0 $X=-550 $Y=-110
X11 1 M1_PO_CDNS_764888589649 $T=-450 1890 0 0 $X=-550 $Y=1770
X12 3 M1_PO_CDNS_764888589649 $T=-40 -2140 0 0 $X=-140 $Y=-2260
X13 1 M1_PO_CDNS_764888589649 $T=-40 1890 0 0 $X=-140 $Y=1770
X14 6 M1_PO_CDNS_764888589649 $T=850 -980 0 0 $X=750 $Y=-1100
X15 5 6 1 5 4 2 pmos1v_CDNS_764888589640 $T=-500 230 0 0 $X=-920 $Y=30
X16 1 5 6 1 4 2 pmos1v_CDNS_764888589640 $T=800 230 0 0 $X=380 $Y=30
X17 5 6 3 5 4 nmos1v_CDNS_764888589641 $T=-500 -1920 0 0 $X=-920 $Y=-2120
X18 3 5 6 3 4 nmos1v_CDNS_764888589641 $T=800 -1920 0 0 $X=380 $Y=-2120
X19 1 2 3 4 inv $T=-1740 -400 0 0 $X=-2220 $Y=-2560
M0 5 1 6 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=-90 $Y=230 $dt=1
M1 5 6 1 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=800 $Y=230 $dt=1
M2 1 6 5 2 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=1210 $Y=230 $dt=1
.ends xor

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764888589642                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764888589642 1 2 3 4 5 6 7 8 9
** N=9 EP=9 FDC=4
M0 2 3 1 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 fw=3.6e-07 sa=1.4e-07 sb=7.55e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=0 $Y=0 $dt=0
M1 4 6 2 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=3.45e-07 sb=5.5e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=410 $Y=0 $dt=0
M2 5 7 4 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.76e-14 AS=5.76e-14 PD=1.04e-06 PS=1.04e-06 fw=3.6e-07 sa=5.5e-07 sb=3.45e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=820 $Y=0 $dt=0
M3 8 9 5 4 g45n1svt L=4.5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 fw=3.6e-07 sa=7.55e-07 sb=1.4e-07 sca=4.15332 scb=0.000375834 scc=2.03107e-07 $X=1230 $Y=0 $dt=0
.ends nmos1v_CDNS_764888589642

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764888589643                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764888589643 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=4
M0 2 4 1 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=7.55e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=0 $Y=0 $dt=1
M1 3 5 2 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=5.5e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=410 $Y=0 $dt=1
M2 6 8 3 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.152e-13 PD=1.76e-06 PS=1.76e-06 fw=7.2e-07 sa=5.5e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=820 $Y=0 $dt=1
M3 7 9 6 11 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=7.55e-07 sb=1.4e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=1230 $Y=0 $dt=1
.ends pmos1v_CDNS_764888589643

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: fa_co_network                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt fa_co_network 1 2 3 4 5 6 7 8 9 10
+ 11
** N=11 EP=11 FDC=8
X0 1 M2_M1_CDNS_764888589643 $T=-830 -970 0 0 $X=-910 $Y=-1100
X1 2 M2_M1_CDNS_764888589643 $T=-220 -60 0 0 $X=-300 $Y=-190
X2 2 M2_M1_CDNS_764888589643 $T=200 730 0 0 $X=120 $Y=600
X3 1 M2_M1_CDNS_764888589643 $T=810 -970 0 0 $X=730 $Y=-1100
X4 2 M1_PO_CDNS_764888589649 $T=-220 -60 0 0 $X=-320 $Y=-180
X5 5 M1_PO_CDNS_764888589649 $T=-210 730 0 0 $X=-310 $Y=610
X6 5 M1_PO_CDNS_764888589649 $T=190 -60 0 0 $X=90 $Y=-180
X7 2 M1_PO_CDNS_764888589649 $T=200 730 0 0 $X=100 $Y=610
X8 4 M1_NWELL_CDNS_7648885896412 $T=-10 2990 0 0 $X=-430 $Y=2690
X9 3 M1_PO_CDNS_7648885896413 $T=-590 550 0 0 $X=-690 $Y=190
X10 7 M1_PO_CDNS_7648885896413 $T=570 550 0 0 $X=470 $Y=190
X11 6 M1_PSUB_CDNS_7648885896414 $T=0 -1600 0 0 $X=-380 $Y=-1740
X12 1 8 3 6 9 2 5 1 7 nmos1v_CDNS_764888589642 $T=-670 -1100 0 0 $X=-1090 $Y=-1300
X13 1 10 4 3 5 11 1 2 7 6
+ 4 pmos1v_CDNS_764888589643 $T=-670 1050 0 0 $X=-1090 $Y=850
.ends fa_co_network

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder_auto                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder_auto 3 7 2 6 8 1 10
** N=15 EP=7 FDC=36
X0 1 M2_M1_CDNS_764888589640 $T=7490 13680 0 0 $X=7360 $Y=13550
X1 2 M2_M1_CDNS_764888589640 $T=8640 11120 0 0 $X=8510 $Y=10990
X2 2 M2_M1_CDNS_764888589640 $T=11340 11400 0 0 $X=11210 $Y=11270
X3 1 M2_M1_CDNS_764888589641 $T=4440 13680 0 0 $X=4310 $Y=13550
X4 2 M3_M2_CDNS_764888589642 $T=8320 11120 0 0 $X=8190 $Y=10990
X5 2 M3_M2_CDNS_764888589642 $T=11130 11400 0 0 $X=11000 $Y=11270
X6 3 M2_M1_CDNS_764888589643 $T=6270 10830 0 0 $X=6190 $Y=10700
X7 4 M2_M1_CDNS_764888589643 $T=10550 10140 0 0 $X=10470 $Y=10010
X8 5 M2_M1_CDNS_764888589643 $T=10550 12850 0 0 $X=10470 $Y=12720
X9 1 M2_M1_CDNS_764888589643 $T=11840 13730 0 0 $X=11760 $Y=13600
X10 4 M2_M1_CDNS_764888589643 $T=12060 10700 0 0 $X=11980 $Y=10570
X11 3 M2_M1_CDNS_764888589643 $T=12410 11080 0 0 $X=12330 $Y=10950
X12 6 M2_M1_CDNS_764888589643 $T=13940 11270 0 0 $X=13860 $Y=11140
X13 7 M3_M2_CDNS_764888589644 $T=3290 11620 0 0 $X=3210 $Y=11490
X14 3 M3_M2_CDNS_764888589644 $T=6810 10840 0 0 $X=6730 $Y=10710
X15 8 M3_M2_CDNS_764888589644 $T=10140 12520 0 0 $X=10060 $Y=12390
X16 3 M3_M2_CDNS_764888589644 $T=12430 10700 0 0 $X=12350 $Y=10570
X17 6 M3_M2_CDNS_764888589644 $T=13940 11270 0 0 $X=13860 $Y=11140
X18 3 M4_M3_CDNS_764888589645 $T=8000 10840 0 0 $X=7920 $Y=10710
X19 3 M4_M3_CDNS_764888589645 $T=11160 10730 0 0 $X=11080 $Y=10600
X20 9 1 6 10 inv $T=13370 11170 0 0 $X=12890 $Y=9010
X21 7 1 11 10 5 3 xor $T=5190 11570 0 0 $X=2970 $Y=9010
X22 5 1 4 10 8 2 xor $T=9090 11570 0 0 $X=6870 $Y=9010
X23 9 5 2 1 4 10 3 12 13 14
+ 15 fa_co_network $T=11860 10750 0 0 $X=10770 $Y=9010
M0 11 7 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=3390 $Y=11800 $dt=1
M1 1 7 11 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=3800 $Y=11800 $dt=1
M2 3 7 5 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.8711 scb=0.0135953 scc=0.00231129 $X=4690 $Y=11800 $dt=1
M3 4 5 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7290 $Y=11800 $dt=1
M4 1 5 4 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=7700 $Y=11800 $dt=1
M5 2 5 8 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=25.5135 scb=0.01349 scc=0.00231127 $X=8590 $Y=11800 $dt=1
M6 6 9 1 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.152e-13 AS=1.008e-13 PD=1.76e-06 PS=1.72e-06 fw=7.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.0436 scb=0.0194268 scc=0.00239616 $X=13310 $Y=11800 $dt=1
M7 1 9 6 1 g45p1svt L=4.5e-08 W=7.2e-07 AD=1.008e-13 AS=1.152e-13 PD=1.72e-06 PS=1.76e-06 fw=7.2e-07 sa=3.45e-07 sb=1.4e-07 sca=44.9648 scb=0.0375178 scc=0.00495812 $X=13720 $Y=11800 $dt=1
.ends full_adder_auto
